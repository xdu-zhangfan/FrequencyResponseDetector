// Verilog netlist created by Tang Dynasty v5.6.71036
// Mon Jul 10 11:12:22 2023

`timescale 1ns / 1ps
module dds_phy
  (
  clk,
  fword,
  pword,
  rst_n,
  phase_out,
  rdy,
  wave_cos,
  wave_sin
  );

  input clk;
  input [31:0] fword;
  input [31:0] pword;
  input rst_n;
  output [31:0] phase_out;
  output rdy;
  output [13:0] wave_cos;
  output [13:0] wave_sin;

  parameter FREC_OUT = 1000000;
  parameter FREC_SYS = 120000000;
  parameter LENTH_ROM = 4096;
  parameter W_DOUT = 14;
  parameter W_PHASE = 32;
  parameter W_PHASE_ANGLE = 14;
  // localparam PHA_INC = 35791394;
  // localparam W_JITTER = 2;
  wire [31:0] al_4c12045b;
  wire [31:0] al_7521c31;
  wire [10:0] al_80d2564a;
  wire [10:0] al_35c5bf4a;
  wire [10:0] al_b33e7450;
  wire [10:0] al_8aaaf100;
  wire [10:0] al_6790cfef;
  wire [10:0] al_8378b540;
  wire [12:0] al_7cb3139;
  wire [12:0] al_defcae67;
  wire [12:0] al_582c7f1a;
  wire [11:0] al_fcd55aa0;
  wire [12:0] al_75776e99;
  wire [12:0] al_e1c1520b;
  wire [12:0] al_7c6da17f;
  wire [11:0] al_d0d95c2b;
  wire [31:0] al_5e800bf9;
  wire [31:0] al_2adbf503;
  wire [31:0] al_ac33d53a;
  wire [31:0] al_1ca72219;
  wire [31:0] al_8fc74dd1;
  wire [11:0] al_50d27df2;
  wire [13:0] al_3bc6703c;
  wire [31:0] al_45f60c58;
  wire [11:0] al_a07945e6;
  wire [11:0] al_ef10e9eb;
  wire [31:0] al_bf05573;
  wire [11:0] al_bf62f43;
  wire [11:0] al_1db9833e;
  wire [11:0] al_aeba03f9;
  wire [31:0] al_b84f9223;
  wire [11:0] al_2c65e87;
  wire [11:0] al_9644e37b;
  wire [31:0] al_8fd1686;
  wire [11:0] al_ff8d588f;
  wire [11:0] al_b0376e91;
  wire [31:0] al_4fdd6779;
  wire [11:0] al_e765e4ce;
  wire [31:0] al_411d7869;
  wire [31:0] al_347def8c;
  wire [31:0] al_2fc0f064;
  wire [13:0] al_6b994b8c;
  wire [31:0] al_cc82cb7d;
  wire [13:0] al_bc5c8fc3;
  wire [31:0] al_747bea5;
  wire al_eabcde5c;
  wire al_c129e0ce;
  wire al_a91ea309;
  wire al_60d44b4;
  wire al_e3ba0d71;
  wire al_fe0dc866;
  wire al_d034bb7c;
  wire al_59f8c17e;
  wire al_956f61e8;
  wire al_9683e9e9;
  wire al_de15ce6c;
  wire al_bc99628c;
  wire al_646ebcc2;
  wire al_85a14d9;
  wire al_3062c0e5;
  wire al_4cd31cc3;
  wire al_7ac21880;
  wire al_f522446b;
  wire al_90e0f7f4;
  wire al_794cef0c;
  wire al_8b35208e;
  wire al_7fb0038c;
  wire al_e3688d46;
  wire al_ac0ba0da;
  wire al_48f8b31c;
  wire al_85c6bbf1;
  wire al_df2b9fd;
  wire al_8b37f3ea;
  wire al_681a20da;
  wire al_7ee6fbef;
  wire al_bc7eb654;
  wire al_2c954a69;
  wire al_b898adc0;
  wire al_48222c42;
  wire al_ac0e8578;
  wire al_71a81d55;
  wire al_eb089a18;
  wire al_d12b8278;
  wire al_2abb4e54;
  wire al_1d87f1e2;
  wire al_6b7ab472;
  wire al_a5d9ceb0;
  wire al_39b072a6;
  wire al_6d449e6d;
  wire al_e4e44f79;
  wire al_1cf3a40d;
  wire al_aa070a2;
  wire al_5e40219b;
  wire al_4c3de7a8;
  wire al_554d4691;
  wire al_d1a163c3;
  wire al_dcd96e0b;
  wire al_50010de7;
  wire al_3d64a0b5;
  wire al_e497746;
  wire al_dafddd54;
  wire al_b52f0f62;
  wire al_211ae938;
  wire al_395d66fa;
  wire al_a5a39f01;
  wire al_29a49a6c;
  wire al_92bb71b8;
  wire al_71e1cc55;
  wire al_31c20af0;
  wire al_dc38bdb4;
  wire al_76e04b4c;
  wire al_cb080167;
  wire al_b00ea7b0;
  wire al_dac79980;
  wire al_cffcd924;
  wire al_51ee9de4;
  wire al_17cd6e3d;
  wire al_7f59913d;
  wire al_7b778bed;
  wire al_3863a70c;
  wire al_5d0f242;
  wire al_fdfe386c;
  wire al_a206a928;
  wire al_2e229782;
  wire al_6096bb6;
  wire al_8dec1170;
  wire al_31cdbd57;
  wire al_c667bd4e;
  wire al_4252b029;
  wire al_b3cdd3bf;
  wire al_e5086b32;
  wire al_85b84194;
  wire al_697e49b8;
  wire al_a7bae841;
  wire al_a41fb992;
  wire al_7c9c9a92;
  wire al_c67d742d;
  wire al_d8746be;
  wire al_157c7876;
  wire al_ee0853c4;
  wire al_7d7c5bcf;
  wire al_76b376c0;
  wire al_42b3f135;
  wire al_dee438f1;
  wire al_f2f78b17;
  wire al_6793a1ac;
  wire al_8ff3cabd;
  wire al_d61e6baf;
  wire al_6c03ab68;
  wire al_4714f41a;
  wire al_8d0c9e0b;
  wire al_fefa949f;
  wire al_ef086a54;
  wire al_8f38553e;
  wire al_85982818;
  wire al_3c9ea8d3;
  wire al_38c1801c;
  wire al_988c595c;
  wire al_e0f22df3;
  wire al_2eab2555;
  wire al_ae82e036;
  wire al_408f5b70;
  wire al_3fc95884;
  wire al_68d1991b;
  wire al_502834ef;
  wire al_5f378f79;
  wire al_8b83adde;
  wire al_fe665c1c;
  wire al_facfca0b;
  wire al_ee9aabaa;
  wire al_9ec1c974;
  wire al_bae62995;
  wire al_72d4aeb7;
  wire al_16154cc8;
  wire al_c8187df2;
  wire al_2866f959;
  wire al_6d9cf46e;
  wire al_8d3c91f3;
  wire al_124cb870;
  wire al_1aefe382;
  wire al_63190405;
  wire al_25fbcbb5;
  wire al_8e2f713c;
  wire al_5fbe7497;

  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_45d6eb2b (
    .a(1'b0),
    .o({al_d61e6baf,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed0aa007 (
    .a(1'b0),
    .b(al_7cb3139[0]),
    .c(al_d61e6baf),
    .o({al_6c03ab68,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b71aa3e2 (
    .a(1'b0),
    .b(al_7cb3139[1]),
    .c(al_6c03ab68),
    .o({al_4714f41a,al_cc82cb7d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59450c7f (
    .a(1'b0),
    .b(al_7cb3139[2]),
    .c(al_4714f41a),
    .o({al_8d0c9e0b,al_cc82cb7d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c728b2ea (
    .a(1'b0),
    .b(al_7cb3139[3]),
    .c(al_8d0c9e0b),
    .o({al_fefa949f,al_cc82cb7d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_71a9d773 (
    .a(1'b0),
    .b(al_7cb3139[4]),
    .c(al_fefa949f),
    .o({al_ef086a54,al_cc82cb7d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_34dc8e91 (
    .a(1'b0),
    .b(al_7cb3139[5]),
    .c(al_ef086a54),
    .o({al_8f38553e,al_cc82cb7d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b58d2e52 (
    .a(1'b0),
    .b(al_7cb3139[6]),
    .c(al_8f38553e),
    .o({al_85982818,al_cc82cb7d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d200bc7 (
    .a(1'b0),
    .b(al_7cb3139[7]),
    .c(al_85982818),
    .o({al_3c9ea8d3,al_cc82cb7d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b8bdd9 (
    .a(1'b0),
    .b(al_7cb3139[8]),
    .c(al_3c9ea8d3),
    .o({al_38c1801c,al_cc82cb7d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d9d9d7a (
    .a(1'b0),
    .b(al_7cb3139[9]),
    .c(al_38c1801c),
    .o({al_988c595c,al_cc82cb7d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9cce3cfb (
    .a(1'b0),
    .b(al_7cb3139[10]),
    .c(al_988c595c),
    .o({al_e0f22df3,al_cc82cb7d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55e53dc7 (
    .a(1'b0),
    .b(al_7cb3139[11]),
    .c(al_e0f22df3),
    .o({al_2eab2555,al_cc82cb7d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1305ee25 (
    .a(1'b0),
    .b(al_7cb3139[12]),
    .c(al_2eab2555),
    .o({al_ae82e036,al_cc82cb7d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58d3b56c (
    .c(al_ae82e036),
    .o({open_n6,al_cc82cb7d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1eb6e7f4 (
    .a(1'b0),
    .o({al_408f5b70,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5070be8a (
    .a(1'b0),
    .b(al_8fc74dd1[18]),
    .c(al_408f5b70),
    .o({al_3fc95884,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_199b9a22 (
    .a(1'b0),
    .b(al_8fc74dd1[19]),
    .c(al_3fc95884),
    .o({al_68d1991b,al_3bc6703c[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_194c9640 (
    .a(1'b0),
    .b(al_8fc74dd1[20]),
    .c(al_68d1991b),
    .o({al_502834ef,al_3bc6703c[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fe0a249 (
    .a(1'b0),
    .b(al_8fc74dd1[21]),
    .c(al_502834ef),
    .o({al_5f378f79,al_3bc6703c[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3d75bc27 (
    .a(1'b0),
    .b(al_8fc74dd1[22]),
    .c(al_5f378f79),
    .o({al_8b83adde,al_3bc6703c[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ad639e (
    .a(1'b0),
    .b(al_8fc74dd1[23]),
    .c(al_8b83adde),
    .o({al_fe665c1c,al_3bc6703c[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aede42cd (
    .a(1'b0),
    .b(al_8fc74dd1[24]),
    .c(al_fe665c1c),
    .o({al_facfca0b,al_3bc6703c[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1252e212 (
    .a(1'b0),
    .b(al_8fc74dd1[25]),
    .c(al_facfca0b),
    .o({al_ee9aabaa,al_3bc6703c[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_802d6d3e (
    .a(1'b0),
    .b(al_8fc74dd1[26]),
    .c(al_ee9aabaa),
    .o({al_9ec1c974,al_3bc6703c[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f07c543 (
    .a(1'b0),
    .b(al_8fc74dd1[27]),
    .c(al_9ec1c974),
    .o({al_bae62995,al_3bc6703c[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50fd806a (
    .a(1'b0),
    .b(al_8fc74dd1[28]),
    .c(al_bae62995),
    .o({al_72d4aeb7,al_3bc6703c[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5eea9400 (
    .a(1'b0),
    .b(al_8fc74dd1[29]),
    .c(al_72d4aeb7),
    .o({open_n11,al_3bc6703c[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_8c9c8dcf (
    .a(1'b0),
    .o({al_a7bae841,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7be4e5a6 (
    .a(1'b0),
    .b(al_75776e99[0]),
    .c(al_a7bae841),
    .o({al_a41fb992,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ac6f968 (
    .a(1'b0),
    .b(al_75776e99[1]),
    .c(al_a41fb992),
    .o({al_7c9c9a92,al_747bea5[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_66955c (
    .a(1'b0),
    .b(al_75776e99[2]),
    .c(al_7c9c9a92),
    .o({al_c67d742d,al_747bea5[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_75a95cba (
    .a(1'b0),
    .b(al_75776e99[3]),
    .c(al_c67d742d),
    .o({al_d8746be,al_747bea5[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7019c95 (
    .a(1'b0),
    .b(al_75776e99[4]),
    .c(al_d8746be),
    .o({al_157c7876,al_747bea5[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_510eb9ca (
    .a(1'b0),
    .b(al_75776e99[5]),
    .c(al_157c7876),
    .o({al_ee0853c4,al_747bea5[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aec64ec2 (
    .a(1'b0),
    .b(al_75776e99[6]),
    .c(al_ee0853c4),
    .o({al_7d7c5bcf,al_747bea5[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fe6f5db3 (
    .a(1'b0),
    .b(al_75776e99[7]),
    .c(al_7d7c5bcf),
    .o({al_76b376c0,al_747bea5[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d76ede99 (
    .a(1'b0),
    .b(al_75776e99[8]),
    .c(al_76b376c0),
    .o({al_42b3f135,al_747bea5[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e3b383d9 (
    .a(1'b0),
    .b(al_75776e99[9]),
    .c(al_42b3f135),
    .o({al_dee438f1,al_747bea5[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1bbb11e (
    .a(1'b0),
    .b(al_75776e99[10]),
    .c(al_dee438f1),
    .o({al_f2f78b17,al_747bea5[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a69b355d (
    .a(1'b0),
    .b(al_75776e99[11]),
    .c(al_f2f78b17),
    .o({al_6793a1ac,al_747bea5[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a628ec5e (
    .a(1'b0),
    .b(al_75776e99[12]),
    .c(al_6793a1ac),
    .o({al_8ff3cabd,al_747bea5[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fde77d46 (
    .c(al_8ff3cabd),
    .o({open_n18,al_747bea5[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b22ad72b (
    .a(al_8378b540[8]),
    .b(al_e765e4ce[7]),
    .c(al_59f8c17e),
    .o({al_956f61e8,al_d0d95c2b[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37642c3c (
    .a(al_8378b540[9]),
    .b(al_e765e4ce[8]),
    .c(al_956f61e8),
    .o({al_9683e9e9,al_d0d95c2b[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a06a895b (
    .a(al_8378b540[10]),
    .b(al_e765e4ce[9]),
    .c(al_9683e9e9),
    .o({al_de15ce6c,al_d0d95c2b[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_877fa7f9 (
    .a(1'b0),
    .b(al_e765e4ce[10]),
    .c(al_de15ce6c),
    .o({al_bc99628c,al_d0d95c2b[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2d21f01f (
    .a(1'b0),
    .b(al_e765e4ce[11]),
    .c(al_bc99628c),
    .o({open_n19,al_d0d95c2b[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_41335dfd (
    .a(1'b0),
    .o({al_eabcde5c,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_513090b3 (
    .a(al_8378b540[1]),
    .b(al_b0376e91[0]),
    .c(al_eabcde5c),
    .o({al_c129e0ce,al_d0d95c2b[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6708c65 (
    .a(al_8378b540[2]),
    .b(al_e765e4ce[1]),
    .c(al_c129e0ce),
    .o({al_a91ea309,al_d0d95c2b[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8a72a648 (
    .a(al_8378b540[3]),
    .b(al_e765e4ce[2]),
    .c(al_a91ea309),
    .o({al_60d44b4,al_d0d95c2b[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a4d828f2 (
    .a(al_8378b540[4]),
    .b(al_e765e4ce[3]),
    .c(al_60d44b4),
    .o({al_e3ba0d71,al_d0d95c2b[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8b186716 (
    .a(al_8378b540[5]),
    .b(al_e765e4ce[4]),
    .c(al_e3ba0d71),
    .o({al_fe0dc866,al_d0d95c2b[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3d917c9c (
    .a(al_8378b540[6]),
    .b(al_e765e4ce[5]),
    .c(al_fe0dc866),
    .o({al_d034bb7c,al_d0d95c2b[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e7664728 (
    .a(al_8378b540[7]),
    .b(al_e765e4ce[6]),
    .c(al_d034bb7c),
    .o({al_59f8c17e,al_d0d95c2b[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_447e8c98 (
    .a(1'b0),
    .o({al_646ebcc2,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dfe88b8b (
    .a(al_4c12045b[8]),
    .b(al_5e800bf9[8]),
    .c(al_8b35208e),
    .o({al_7fb0038c,al_7521c31[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_25ea18a5 (
    .a(al_4c12045b[9]),
    .b(al_5e800bf9[9]),
    .c(al_7fb0038c),
    .o({al_e3688d46,al_7521c31[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_102c5891 (
    .a(al_4c12045b[10]),
    .b(al_5e800bf9[10]),
    .c(al_e3688d46),
    .o({al_ac0ba0da,al_7521c31[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cfaa08b6 (
    .a(al_4c12045b[11]),
    .b(al_5e800bf9[11]),
    .c(al_ac0ba0da),
    .o({al_48f8b31c,al_7521c31[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_33d1b43 (
    .a(al_4c12045b[12]),
    .b(al_5e800bf9[12]),
    .c(al_48f8b31c),
    .o({al_85c6bbf1,al_7521c31[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d9268e1f (
    .a(al_4c12045b[13]),
    .b(al_5e800bf9[13]),
    .c(al_85c6bbf1),
    .o({al_df2b9fd,al_7521c31[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8d2d7bf1 (
    .a(al_4c12045b[14]),
    .b(al_5e800bf9[14]),
    .c(al_df2b9fd),
    .o({al_8b37f3ea,al_7521c31[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37795e33 (
    .a(al_4c12045b[15]),
    .b(al_5e800bf9[15]),
    .c(al_8b37f3ea),
    .o({al_681a20da,al_7521c31[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_819cb1a2 (
    .a(al_4c12045b[16]),
    .b(al_5e800bf9[16]),
    .c(al_681a20da),
    .o({al_7ee6fbef,al_7521c31[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6df20a54 (
    .a(al_4c12045b[17]),
    .b(al_5e800bf9[17]),
    .c(al_7ee6fbef),
    .o({al_bc7eb654,al_7521c31[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4cc92009 (
    .a(al_4c12045b[0]),
    .b(al_5e800bf9[0]),
    .c(al_646ebcc2),
    .o({al_85a14d9,al_7521c31[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8d80c396 (
    .a(al_4c12045b[18]),
    .b(al_5e800bf9[18]),
    .c(al_bc7eb654),
    .o({al_2c954a69,al_7521c31[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_22dfbf6 (
    .a(al_4c12045b[19]),
    .b(al_5e800bf9[19]),
    .c(al_2c954a69),
    .o({al_b898adc0,al_7521c31[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b6ce109b (
    .a(al_4c12045b[20]),
    .b(al_5e800bf9[20]),
    .c(al_b898adc0),
    .o({al_48222c42,al_7521c31[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3be7cdd2 (
    .a(al_4c12045b[21]),
    .b(al_5e800bf9[21]),
    .c(al_48222c42),
    .o({al_ac0e8578,al_7521c31[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_abc5c8fc (
    .a(al_4c12045b[22]),
    .b(al_5e800bf9[22]),
    .c(al_ac0e8578),
    .o({al_71a81d55,al_7521c31[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_35dee330 (
    .a(al_4c12045b[23]),
    .b(al_5e800bf9[23]),
    .c(al_71a81d55),
    .o({al_eb089a18,al_7521c31[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6a3e0a0 (
    .a(al_4c12045b[24]),
    .b(al_5e800bf9[24]),
    .c(al_eb089a18),
    .o({al_d12b8278,al_7521c31[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cea749b0 (
    .a(al_4c12045b[25]),
    .b(al_5e800bf9[25]),
    .c(al_d12b8278),
    .o({al_2abb4e54,al_7521c31[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6d66ee19 (
    .a(al_4c12045b[26]),
    .b(al_5e800bf9[26]),
    .c(al_2abb4e54),
    .o({al_1d87f1e2,al_7521c31[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3bbe2c91 (
    .a(al_4c12045b[27]),
    .b(al_5e800bf9[27]),
    .c(al_1d87f1e2),
    .o({al_6b7ab472,al_7521c31[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b3abc203 (
    .a(al_4c12045b[1]),
    .b(al_5e800bf9[1]),
    .c(al_85a14d9),
    .o({al_3062c0e5,al_7521c31[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_41d36f2b (
    .a(al_4c12045b[28]),
    .b(al_5e800bf9[28]),
    .c(al_6b7ab472),
    .o({al_a5d9ceb0,al_7521c31[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8b54afaf (
    .a(al_4c12045b[29]),
    .b(al_5e800bf9[29]),
    .c(al_a5d9ceb0),
    .o({al_39b072a6,al_7521c31[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_90b1a19d (
    .a(al_4c12045b[30]),
    .b(al_5e800bf9[30]),
    .c(al_39b072a6),
    .o({al_6d449e6d,al_7521c31[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e56607bb (
    .a(al_4c12045b[31]),
    .b(al_5e800bf9[31]),
    .c(al_6d449e6d),
    .o({open_n26,al_7521c31[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9a29b387 (
    .a(al_4c12045b[2]),
    .b(al_5e800bf9[2]),
    .c(al_3062c0e5),
    .o({al_4cd31cc3,al_7521c31[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f8409470 (
    .a(al_4c12045b[3]),
    .b(al_5e800bf9[3]),
    .c(al_4cd31cc3),
    .o({al_7ac21880,al_7521c31[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_68cc8618 (
    .a(al_4c12045b[4]),
    .b(al_5e800bf9[4]),
    .c(al_7ac21880),
    .o({al_f522446b,al_7521c31[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7669cd7d (
    .a(al_4c12045b[5]),
    .b(al_5e800bf9[5]),
    .c(al_f522446b),
    .o({al_90e0f7f4,al_7521c31[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7b766b13 (
    .a(al_4c12045b[6]),
    .b(al_5e800bf9[6]),
    .c(al_90e0f7f4),
    .o({al_794cef0c,al_7521c31[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dac99e8a (
    .a(al_4c12045b[7]),
    .b(al_5e800bf9[7]),
    .c(al_794cef0c),
    .o({al_8b35208e,al_7521c31[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c22ee456 (
    .a(al_b33e7450[8]),
    .b(al_b0376e91[7]),
    .c(al_dcd96e0b),
    .o({al_50010de7,al_fcd55aa0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4f8c6b2 (
    .a(al_b33e7450[9]),
    .b(al_b0376e91[8]),
    .c(al_50010de7),
    .o({al_3d64a0b5,al_fcd55aa0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_251c9501 (
    .a(al_b33e7450[10]),
    .b(al_b0376e91[9]),
    .c(al_3d64a0b5),
    .o({al_e497746,al_fcd55aa0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b10f851 (
    .a(1'b0),
    .b(al_b0376e91[10]),
    .c(al_e497746),
    .o({al_dafddd54,al_fcd55aa0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f6074d25 (
    .a(1'b0),
    .b(al_b0376e91[11]),
    .c(al_dafddd54),
    .o({open_n27,al_fcd55aa0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_542d5c78 (
    .a(1'b0),
    .o({al_e4e44f79,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a685a1be (
    .a(al_b33e7450[1]),
    .b(al_b0376e91[0]),
    .c(al_e4e44f79),
    .o({al_1cf3a40d,al_fcd55aa0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cda14380 (
    .a(al_b33e7450[2]),
    .b(al_b0376e91[1]),
    .c(al_1cf3a40d),
    .o({al_aa070a2,al_fcd55aa0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f54c3dbb (
    .a(al_b33e7450[3]),
    .b(al_b0376e91[2]),
    .c(al_aa070a2),
    .o({al_5e40219b,al_fcd55aa0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c9b145c3 (
    .a(al_b33e7450[4]),
    .b(al_b0376e91[3]),
    .c(al_5e40219b),
    .o({al_4c3de7a8,al_fcd55aa0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_85743617 (
    .a(al_b33e7450[5]),
    .b(al_b0376e91[4]),
    .c(al_4c3de7a8),
    .o({al_554d4691,al_fcd55aa0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ad670f93 (
    .a(al_b33e7450[6]),
    .b(al_b0376e91[5]),
    .c(al_554d4691),
    .o({al_d1a163c3,al_fcd55aa0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec16458c (
    .a(al_b33e7450[7]),
    .b(al_b0376e91[6]),
    .c(al_d1a163c3),
    .o({al_dcd96e0b,al_fcd55aa0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_1e2e84c8 (
    .a(1'b0),
    .o({al_b52f0f62,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9741ddb6 (
    .a(al_4c12045b[8]),
    .b(al_2fc0f064[8]),
    .c(al_dc38bdb4),
    .o({al_76e04b4c,al_ac33d53a[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cb2d7da6 (
    .a(al_4c12045b[9]),
    .b(al_2fc0f064[9]),
    .c(al_76e04b4c),
    .o({al_cb080167,al_ac33d53a[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a5d95d17 (
    .a(al_4c12045b[10]),
    .b(al_2fc0f064[10]),
    .c(al_cb080167),
    .o({al_b00ea7b0,al_ac33d53a[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c7cc56f4 (
    .a(al_4c12045b[11]),
    .b(al_2fc0f064[11]),
    .c(al_b00ea7b0),
    .o({al_dac79980,al_ac33d53a[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_65bf2a28 (
    .a(al_4c12045b[12]),
    .b(al_2fc0f064[12]),
    .c(al_dac79980),
    .o({al_cffcd924,al_ac33d53a[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c4008c1d (
    .a(al_4c12045b[13]),
    .b(al_2fc0f064[13]),
    .c(al_cffcd924),
    .o({al_51ee9de4,al_ac33d53a[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_66a06386 (
    .a(al_4c12045b[14]),
    .b(al_2fc0f064[14]),
    .c(al_51ee9de4),
    .o({al_17cd6e3d,al_ac33d53a[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6e1f94b1 (
    .a(al_4c12045b[15]),
    .b(al_2fc0f064[15]),
    .c(al_17cd6e3d),
    .o({al_7f59913d,al_ac33d53a[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e6d64658 (
    .a(al_4c12045b[16]),
    .b(al_2fc0f064[16]),
    .c(al_7f59913d),
    .o({al_7b778bed,al_ac33d53a[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9266bf3 (
    .a(al_4c12045b[17]),
    .b(al_2fc0f064[17]),
    .c(al_7b778bed),
    .o({al_3863a70c,al_ac33d53a[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c0083060 (
    .a(al_4c12045b[0]),
    .b(al_2fc0f064[0]),
    .c(al_b52f0f62),
    .o({al_211ae938,al_ac33d53a[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3ee46d9 (
    .a(al_4c12045b[18]),
    .b(al_2fc0f064[18]),
    .c(al_3863a70c),
    .o({al_5d0f242,al_ac33d53a[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9cba80ba (
    .a(al_4c12045b[19]),
    .b(al_2fc0f064[19]),
    .c(al_5d0f242),
    .o({al_fdfe386c,al_ac33d53a[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_77660ab8 (
    .a(al_4c12045b[20]),
    .b(al_2fc0f064[20]),
    .c(al_fdfe386c),
    .o({al_a206a928,al_ac33d53a[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1783073b (
    .a(al_4c12045b[21]),
    .b(al_2fc0f064[21]),
    .c(al_a206a928),
    .o({al_2e229782,al_ac33d53a[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2b31b946 (
    .a(al_4c12045b[22]),
    .b(al_2fc0f064[22]),
    .c(al_2e229782),
    .o({al_6096bb6,al_ac33d53a[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_caf49207 (
    .a(al_4c12045b[23]),
    .b(al_2fc0f064[23]),
    .c(al_6096bb6),
    .o({al_8dec1170,al_ac33d53a[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b654913e (
    .a(al_4c12045b[24]),
    .b(al_2fc0f064[24]),
    .c(al_8dec1170),
    .o({al_31cdbd57,al_ac33d53a[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_995b24e9 (
    .a(al_4c12045b[25]),
    .b(al_2fc0f064[25]),
    .c(al_31cdbd57),
    .o({al_c667bd4e,al_ac33d53a[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_32cbfc52 (
    .a(al_4c12045b[26]),
    .b(al_2fc0f064[26]),
    .c(al_c667bd4e),
    .o({al_4252b029,al_ac33d53a[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b0617d4d (
    .a(al_4c12045b[27]),
    .b(al_2fc0f064[27]),
    .c(al_4252b029),
    .o({al_b3cdd3bf,al_ac33d53a[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f174f118 (
    .a(al_4c12045b[1]),
    .b(al_2fc0f064[1]),
    .c(al_211ae938),
    .o({al_395d66fa,al_ac33d53a[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ac9f8517 (
    .a(al_4c12045b[28]),
    .b(al_2fc0f064[28]),
    .c(al_b3cdd3bf),
    .o({al_e5086b32,al_ac33d53a[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9a75dbc (
    .a(al_4c12045b[29]),
    .b(al_2fc0f064[29]),
    .c(al_e5086b32),
    .o({al_85b84194,al_ac33d53a[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bd641f50 (
    .a(al_4c12045b[30]),
    .b(al_2fc0f064[30]),
    .c(al_85b84194),
    .o({al_697e49b8,al_ac33d53a[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_69967d4f (
    .a(al_4c12045b[31]),
    .b(al_2fc0f064[31]),
    .c(al_697e49b8),
    .o({open_n34,al_ac33d53a[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_65a345c7 (
    .a(al_4c12045b[2]),
    .b(al_2fc0f064[2]),
    .c(al_395d66fa),
    .o({al_a5a39f01,al_ac33d53a[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9fdf7958 (
    .a(al_4c12045b[3]),
    .b(al_2fc0f064[3]),
    .c(al_a5a39f01),
    .o({al_29a49a6c,al_ac33d53a[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cfa89020 (
    .a(al_4c12045b[4]),
    .b(al_2fc0f064[4]),
    .c(al_29a49a6c),
    .o({al_92bb71b8,al_ac33d53a[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d93f603c (
    .a(al_4c12045b[5]),
    .b(al_2fc0f064[5]),
    .c(al_92bb71b8),
    .o({al_71e1cc55,al_ac33d53a[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_407e6c0 (
    .a(al_4c12045b[6]),
    .b(al_2fc0f064[6]),
    .c(al_71e1cc55),
    .o({al_31c20af0,al_ac33d53a[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8c5662f0 (
    .a(al_4c12045b[7]),
    .b(al_2fc0f064[7]),
    .c(al_31c20af0),
    .o({al_dc38bdb4,al_ac33d53a[7]}));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_b6dda1b6 (
    .a(al_16154cc8),
    .b(al_582c7f1a[0]),
    .o(al_defcae67[0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_4f679765 (
    .a(al_16154cc8),
    .b(al_582c7f1a[10]),
    .o(al_defcae67[10]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_48e066c2 (
    .a(al_16154cc8),
    .b(al_582c7f1a[11]),
    .o(al_defcae67[11]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_2dfc7b51 (
    .a(al_16154cc8),
    .b(al_582c7f1a[12]),
    .o(al_defcae67[12]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_185bde12 (
    .a(al_16154cc8),
    .b(al_582c7f1a[1]),
    .o(al_defcae67[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_c1988ea (
    .a(al_16154cc8),
    .b(al_582c7f1a[2]),
    .o(al_defcae67[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_3376e1cf (
    .a(al_16154cc8),
    .b(al_582c7f1a[3]),
    .o(al_defcae67[3]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_7c92ce6b (
    .a(al_16154cc8),
    .b(al_582c7f1a[4]),
    .o(al_defcae67[4]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_c465e73f (
    .a(al_16154cc8),
    .b(al_582c7f1a[5]),
    .o(al_defcae67[5]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_41cfedf7 (
    .a(al_16154cc8),
    .b(al_582c7f1a[6]),
    .o(al_defcae67[6]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_253a7f75 (
    .a(al_16154cc8),
    .b(al_582c7f1a[7]),
    .o(al_defcae67[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_f204fdb3 (
    .a(al_16154cc8),
    .b(al_582c7f1a[8]),
    .o(al_defcae67[8]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_2ed468ce (
    .a(al_16154cc8),
    .b(al_582c7f1a[9]),
    .o(al_defcae67[9]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_e7719e5c (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[0]),
    .o(al_e1c1520b[0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_d515b802 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[10]),
    .o(al_e1c1520b[10]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_5da96408 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[11]),
    .o(al_e1c1520b[11]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_60fb8447 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[12]),
    .o(al_e1c1520b[12]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_94a75fe2 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[1]),
    .o(al_e1c1520b[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_b4d9aa1c (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[2]),
    .o(al_e1c1520b[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_9068d8fe (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[3]),
    .o(al_e1c1520b[3]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_4349e479 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[4]),
    .o(al_e1c1520b[4]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_ad9414d2 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[5]),
    .o(al_e1c1520b[5]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_7b95c4a (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[6]),
    .o(al_e1c1520b[6]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_70d41bf2 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[7]),
    .o(al_e1c1520b[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_76e1ae5b (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[8]),
    .o(al_e1c1520b[8]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_f4b7a93 (
    .a(al_8d3c91f3),
    .b(al_7c6da17f[9]),
    .o(al_e1c1520b[9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d525a5fc (
    .a(al_50d27df2[10]),
    .b(al_45f60c58[28]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cc31806d (
    .a(al_50d27df2[11]),
    .b(al_45f60c58[29]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3ca92187 (
    .a(al_50d27df2[1]),
    .b(al_45f60c58[19]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6c1f08da (
    .a(al_50d27df2[2]),
    .b(al_45f60c58[20]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_97b9fe7d (
    .a(al_50d27df2[3]),
    .b(al_45f60c58[21]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2076ca4d (
    .a(al_50d27df2[4]),
    .b(al_45f60c58[22]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_922d1e28 (
    .a(al_50d27df2[5]),
    .b(al_45f60c58[23]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d94f09f6 (
    .a(al_50d27df2[6]),
    .b(al_45f60c58[24]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5004aa34 (
    .a(al_50d27df2[7]),
    .b(al_45f60c58[25]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e444e8da (
    .a(al_50d27df2[8]),
    .b(al_45f60c58[26]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_910a532e (
    .a(al_50d27df2[9]),
    .b(al_45f60c58[27]),
    .c(al_45f60c58[30]),
    .o(al_ef10e9eb[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_641ca39f (
    .a(al_50d27df2[10]),
    .b(al_45f60c58[28]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b93ff035 (
    .a(al_50d27df2[11]),
    .b(al_45f60c58[29]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_408a3a (
    .a(al_50d27df2[1]),
    .b(al_45f60c58[19]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_5d459b87 (
    .a(al_50d27df2[2]),
    .b(al_45f60c58[20]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ffa9fd0d (
    .a(al_50d27df2[3]),
    .b(al_45f60c58[21]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_1323da91 (
    .a(al_50d27df2[4]),
    .b(al_45f60c58[22]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_ee689b0c (
    .a(al_50d27df2[5]),
    .b(al_45f60c58[23]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_46644e49 (
    .a(al_50d27df2[6]),
    .b(al_45f60c58[24]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4a6cd7e0 (
    .a(al_50d27df2[7]),
    .b(al_45f60c58[25]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e18c3a84 (
    .a(al_50d27df2[8]),
    .b(al_45f60c58[26]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_4a0f6d3d (
    .a(al_50d27df2[9]),
    .b(al_45f60c58[27]),
    .c(al_45f60c58[30]),
    .o(al_1db9833e[9]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_e4e62d3e (
    .a(al_b0376e91[0]),
    .b(al_b0376e91[1]),
    .c(al_b0376e91[2]),
    .d(al_b0376e91[3]),
    .e(al_b0376e91[4]),
    .f(al_b0376e91[5]),
    .o(al_2866f959));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_1a563ec2 (
    .a(al_b0376e91[6]),
    .b(al_b0376e91[7]),
    .c(al_b0376e91[8]),
    .d(al_b0376e91[9]),
    .o(al_6d9cf46e));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_7dd8fcfc (
    .a(al_2866f959),
    .b(al_6d9cf46e),
    .c(al_b0376e91[10]),
    .d(al_b0376e91[11]),
    .e(al_4fdd6779[30]),
    .o(al_c8187df2));
  AL_DFF_X al_470a2ab8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_c8187df2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16154cc8));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*~A)"),
    .INIT(64'h0000000000000004))
    al_da3205d2 (
    .a(al_b0376e91[0]),
    .b(al_4fdd6779[30]),
    .c(al_e765e4ce[1]),
    .d(al_e765e4ce[2]),
    .e(al_e765e4ce[3]),
    .f(al_e765e4ce[4]),
    .o(al_1aefe382));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_32865808 (
    .a(al_e765e4ce[5]),
    .b(al_e765e4ce[6]),
    .c(al_e765e4ce[7]),
    .d(al_e765e4ce[8]),
    .o(al_63190405));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_c718c02a (
    .a(al_1aefe382),
    .b(al_63190405),
    .c(al_e765e4ce[9]),
    .d(al_e765e4ce[10]),
    .e(al_e765e4ce[11]),
    .o(al_124cb870));
  AL_DFF_X al_14fec9f5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_124cb870),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d3c91f3));
  PH1_LOGIC_ERAM #(
    //.FORCE_KEEP("OFF"),
    .ADDR_WIDTH_A(12),
    .ADDR_WIDTH_B(12),
    .ASYNC_RESET_RELEASE_A("ASYNC"),
    .ASYNC_RESET_RELEASE_B("ASYNC"),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(4096),
    .DATA_DEPTH_B(4096),
    .DATA_WIDTH_A(11),
    .DATA_WIDTH_B(11),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("20K"),
    .INIT_FILE("init_str:00000000000 10000000000 01000000000 11000000000 10100000000 01100000000 11100000000 00010000000 10010000000 01010000000 11010000000 10110000000 01110000000 11110000000 00001000000 10001000000 01001000000 11001000000 10101000000 01101000000 11101000000 00011000000 10011000000 01011000000 11011000000 10111000000 01111000000 11111000000 00000100000 10000100000 01000100000 11000100000 10100100000 01100100000 11100100000 00010100000 10010100000 01010100000 11010100000 10110100000 01110100000 11110100000 00001100000 10001100000 01001100000 11001100000 00101100000 01101100000 11101100000 00011100000 10011100000 01011100000 11011100000 00111100000 01111100000 11111100000 00000010000 10000010000 01000010000 11000010000 00100010000 01100010000 11100010000 00010010000 10010010000 01010010000 11010010000 00110010000 01110010000 11110010000 00001010000 10001010000 01001010000 11001010000 00101010000 01101010000 11101010000 00011010000 10011010000 01011010000 11011010000 00111010000 01111010000 11111010000 00000110000 10000110000 01000110000 11000110000 00100110000 01100110000 11100110000 00010110000 10010110000 01010110000 11010110000 00110110000 10110110000 11110110000 00001110000 10001110000 01001110000 11001110000 00101110000 10101110000 11101110000 00011110000 10011110000 01011110000 11011110000 00111110000 10111110000 11111110000 00000001000 10000001000 01000001000 11000001000 00100001000 10100001000 11100001000 00010001000 10010001000 01010001000 11010001000 00110001000 10110001000 11110001000 00001001000 10001001000 01001001000 11001001000 00101001000 10101001000 01101001000 00011001000 10011001000 01011001000 11011001000 00111001000 10111001000 01111001000 00000101000 10000101000 01000101000 11000101000 00100101000 10100101000 01100101000 00010101000 10010101000 01010101000 11010101000 00110101000 10110101000 01110101000 11110101000 10001101000 01001101000 11001101000 00101101000 10101101000 01101101000 11101101000 10011101000 01011101000 11011101000 00111101000 10111101000 01111101000 11111101000 00000011000 01000011000 11000011000 00100011000 10100011000 01100011000 11100011000 00010011000 01010011000 11010011000 00110011000 10110011000 01110011000 11110011000 00001011000 01001011000 11001011000 00101011000 10101011000 01101011000 11101011000 00011011000 10011011000 11011011000 00111011000 10111011000 01111011000 11111011000 00000111000 10000111000 01000111000 00100111000 10100111000 01100111000 11100111000 00010111000 10010111000 01010111000 00110111000 10110111000 01110111000 11110111000 00001111000 10001111000 01001111000 11001111000 10101111000 01101111000 11101111000 00011111000 10011111000 01011111000 11011111000 10111111000 01111111000 11111111000 00000000100 10000000100 01000000100 11000000100 00100000100 01100000100 11100000100 00010000100 10010000100 01010000100 11010000100 00110000100 10110000100 11110000100 00001000100 10001000100 01001000100 11001000100 00101000100 10101000100 01101000100 00011000100 10011000100 01011000100 11011000100 00111000100 10111000100 01111000100 11111000100 10000100100 01000100100 11000100100 00100100100 10100100100 01100100100 11100100100 00010100100 01010100100 11010100100 00110100100 10110100100 01110100100 11110100100 00001100100 10001100100 11001100100 00101100100 10101100100 01101100100 11101100100 00011100100 10011100100 01011100100 00111100100 10111100100 01111100100 11111100100 00000010100 10000010100 01000010100 11000010100 10100010100 01100010100 11100010100 00010010100 10010010100 01010010100 11010010100 00110010100 01110010100 11110010100 00001010100 10001010100 01001010100 11001010100 00101010100 10101010100 11101010100 00011010100 10011010100 01011010100 11011010100 00111010100 10111010100 01111010100 11111010100 10000110100 01000110100 11000110100 00100110100 10100110100 01100110100 11100110100 00010110100 01010110100 11010110100 00110110100 10110110100 01110110100 11110110100 00001110100 10001110100 01001110100 00101110100 10101110100 01101110100 11101110100 00011110100 10011110100 01011110100 11011110100 10111110100 01111110100 11111110100 00000001100 10000001100 01000001100 11000001100 00100001100 10100001100 11100001100 00010001100 10010001100 01010001100 11010001100 00110001100 10110001100 01110001100 11110001100 10001001100 01001001100 11001001100 00101001100 10101001100 01101001100 11101001100 00011001100 10011001100 11011001100 00111001100 10111001100 01111001100 11111001100 00000101100 10000101100 01000101100 11000101100 10100101100 01100101100 11100101100 00010101100 10010101100 01010101100 11010101100 00110101100 10110101100 11110101100 00001101100 10001101100 01001101100 11001101100 00101101100 10101101100 01101101100 11101101100 10011101100 01011101100 11011101100 00111101100 10111101100 01111101100 11111101100 00000011100 10000011100 01000011100 00100011100 10100011100 01100011100 11100011100 00010011100 10010011100 01010011100 11010011100 00110011100 10110011100 11110011100 00001011100 10001011100 01001011100 11001011100 00101011100 10101011100 01101011100 11101011100 10011011100 01011011100 11011011100 00111011100 10111011100 01111011100 11111011100 00000111100 10000111100 01000111100 00100111100 10100111100 01100111100 11100111100 00010111100 10010111100 01010111100 11010111100 00110111100 10110111100 01110111100 00001111100 10001111100 01001111100 11001111100 00101111100 10101111100 01101111100 11101111100 00011111100 10011111100 11011111100 00111111100 10111111100 01111111100 11111111100 00000000010 10000000010 01000000010 11000000010 00100000010 10100000010 11100000010 00010000010 10010000010 01010000010 11010000010 00110000010 10110000010 01110000010 11110000010 00001000010 10001000010 11001000010 00101000010 10101000010 01101000010 11101000010 00011000010 10011000010 01011000010 11011000010 00111000010 10111000010 11111000010 00000100010 10000100010 01000100010 11000100010 00100100010 10100100010 01100100010 11100100010 00010100010 10010100010 01010100010 00110100010 10110100010 01110100010 11110100010 00001100010 10001100010 01001100010 11001100010 00101100010 10101100010 01101100010 11101100010 10011100010 01011100010 11011100010 00111100010 10111100010 01111100010 11111100010 00000010010 10000010010 01000010010 11000010010 00100010010 01100010010 11100010010 00010010010 10010010010 01010010010 11010010010 00110010010 10110010010 01110010010 11110010010 00001010010 10001010010 01001010010 00101010010 10101010010 01101010010 11101010010 00011010010 10011010010 01011010010 11011010010 00111010010 10111010010 01111010010 11111010010 00000110010 01000110010 11000110010 00100110010 10100110010 01100110010 11100110010 00010110010 10010110010 01010110010 11010110010 00110110010 10110110010 01110110010 11110110010 10001110010 01001110010 11001110010 00101110010 10101110010 01101110010 11101110010 00011110010 10011110010 01011110010 11011110010 00111110010 10111110010 01111110010 11111110010 10000001010 01000001010 11000001010 00100001010 10100001010 01100001010 11100001010 00010001010 10010001010 01010001010 11010001010 00110001010 10110001010 01110001010 11110001010 00001001010 01001001010 11001001010 00101001010 10101001010 01101001010 11101001010 00011001010 10011001010 01011001010 11011001010 00111001010 10111001010 01111001010 11111001010 00000101010 10000101010 01000101010 00100101010 10100101010 01100101010 11100101010 00010101010 10010101010 01010101010 11010101010 00110101010 10110101010 01110101010 11110101010 00001101010 10001101010 01001101010 11001101010 00101101010 10101101010 11101101010 00011101010 10011101010 01011101010 11011101010 00111101010 10111101010 01111101010 11111101010 00000011010 10000011010 01000011010 11000011010 00100011010 10100011010 01100011010 11100011010 00010011010 10010011010 01010011010 11010011010 10110011010 01110011010 11110011010 00001011010 10001011010 01001011010 11001011010 00101011010 10101011010 01101011010 11101011010 00011011010 10011011010 01011011010 11011011010 00111011010 10111011010 01111011010 11111011010 00000111010 10000111010 01000111010 11000111010 00100111010 01100111010 11100111010 00010111010 10010111010 01010111010 11010111010 00110111010 10110111010 01110111010 11110111010 00001111010 10001111010 01001111010 11001111010 00101111010 10101111010 01101111010 11101111010 00011111010 10011111010 01011111010 11011111010 00111111010 10111111010 01111111010 11111111010 00000000110 10000000110 01000000110 00100000110 10100000110 01100000110 11100000110 00010000110 10010000110 01010000110 11010000110 00110000110 10110000110 01110000110 11110000110 00001000110 10001000110 01001000110 11001000110 00101000110 10101000110 01101000110 11101000110 00011000110 10011000110 01011000110 11011000110 00111000110 10111000110 01111000110 11111000110 00000100110 10000100110 01000100110 11000100110 00100100110 10100100110 01100100110 11100100110 00010100110 10010100110 01010100110 11010100110 00110100110 10110100110 01110100110 11110100110 00001100110 10001100110 01001100110 00101100110 10101100110 01101100110 11101100110 00011100110 10011100110 01011100110 11011100110 00111100110 10111100110 01111100110 11111100110 00000010110 10000010110 01000010110 11000010110 00100010110 10100010110 01100010110 11100010110 00010010110 10010010110 01010010110 11010010110 00110010110 10110010110 01110010110 11110010110 00001010110 10001010110 01001010110 11001010110 00101010110 10101010110 01101010110 11101010110 00011010110 10011010110 01011010110 11011010110 00111010110 10111010110 01111010110 11111010110 00000110110 10000110110 01000110110 11000110110 00100110110 10100110110 01100110110 11100110110 00010110110 10010110110 01010110110 11010110110 00110110110 10110110110 01110110110 11110110110 00001110110 10001110110 01001110110 11001110110 00101110110 10101110110 01101110110 11101110110 00011110110 10011110110 01011110110 11011110110 00111110110 10111110110 01111110110 11111110110 00000001110 10000001110 10000001110 01000001110 11000001110 00100001110 10100001110 01100001110 11100001110 00010001110 10010001110 01010001110 11010001110 00110001110 10110001110 01110001110 11110001110 00001001110 10001001110 01001001110 11001001110 00101001110 10101001110 01101001110 11101001110 00011001110 10011001110 01011001110 11011001110 00111001110 10111001110 01111001110 11111001110 00000101110 10000101110 01000101110 11000101110 00100101110 10100101110 01100101110 11100101110 00010101110 10010101110 01010101110 11010101110 00110101110 00110101110 10110101110 01110101110 11110101110 00001101110 10001101110 01001101110 11001101110 00101101110 10101101110 01101101110 11101101110 00011101110 10011101110 01011101110 11011101110 00111101110 10111101110 01111101110 11111101110 00000011110 10000011110 01000011110 11000011110 00100011110 10100011110 01100011110 11100011110 11100011110 00010011110 10010011110 01010011110 11010011110 00110011110 10110011110 01110011110 11110011110 00001011110 10001011110 01001011110 11001011110 00101011110 10101011110 01101011110 11101011110 00011011110 10011011110 01011011110 11011011110 11011011110 00111011110 10111011110 01111011110 11111011110 00000111110 10000111110 01000111110 11000111110 00100111110 10100111110 01100111110 11100111110 00010111110 10010111110 01010111110 11010111110 00110111110 00110111110 10110111110 01110111110 11110111110 00001111110 10001111110 01001111110 11001111110 00101111110 10101111110 01101111110 11101111110 00011111110 10011111110 01011111110 11011111110 00111111110 00111111110 10111111110 01111111110 11111111110 00000000001 10000000001 01000000001 11000000001 00100000001 10100000001 01100000001 11100000001 00010000001 10010000001 10010000001 01010000001 11010000001 00110000001 10110000001 01110000001 11110000001 00001000001 10001000001 01001000001 11001000001 00101000001 10101000001 01101000001 01101000001 11101000001 00011000001 10011000001 01011000001 11011000001 00111000001 10111000001 01111000001 11111000001 00000100001 10000100001 10000100001 01000100001 11000100001 00100100001 10100100001 01100100001 11100100001 00010100001 10010100001 01010100001 11010100001 00110100001 00110100001 10110100001 01110100001 11110100001 00001100001 10001100001 01001100001 11001100001 00101100001 10101100001 01101100001 01101100001 11101100001 00011100001 10011100001 01011100001 11011100001 00111100001 10111100001 01111100001 11111100001 11111100001 00000010001 10000010001 01000010001 11000010001 00100010001 10100010001 01100010001 11100010001 00010010001 00010010001 10010010001 01010010001 11010010001 00110010001 10110010001 01110010001 11110010001 00001010001 10001010001 10001010001 01001010001 11001010001 00101010001 10101010001 01101010001 11101010001 00011010001 10011010001 10011010001 01011010001 11011010001 00111010001 10111010001 01111010001 11111010001 00000110001 10000110001 10000110001 01000110001 11000110001 00100110001 10100110001 01100110001 11100110001 00010110001 00010110001 10010110001 01010110001 11010110001 00110110001 10110110001 01110110001 11110110001 11110110001 00001110001 10001110001 01001110001 11001110001 00101110001 10101110001 01101110001 01101110001 11101110001 00011110001 10011110001 01011110001 11011110001 00111110001 10111110001 10111110001 01111110001 11111110001 00000001001 10000001001 01000001001 11000001001 11000001001 00100001001 10100001001 01100001001 11100001001 00010001001 10010001001 01010001001 01010001001 11010001001 00110001001 10110001001 01110001001 11110001001 00001001001 00001001001 10001001001 01001001001 11001001001 00101001001 10101001001 01101001001 01101001001 11101001001 00011001001 10011001001 01011001001 11011001001 00111001001 00111001001 10111001001 01111001001 11111001001 00000101001 10000101001 10000101001 01000101001 11000101001 00100101001 10100101001 01100101001 11100101001 11100101001 00010101001 10010101001 01010101001 11010101001 00110101001 00110101001 10110101001 01110101001 11110101001 00001101001 10001101001 10001101001 01001101001 11001101001 00101101001 10101101001 01101101001 01101101001 11101101001 00011101001 10011101001 01011101001 11011101001 11011101001 00111101001 10111101001 01111101001 11111101001 00000011001 00000011001 10000011001 01000011001 11000011001 00100011001 10100011001 10100011001 01100011001 11100011001 00010011001 10010011001 01010011001 01010011001 11010011001 00110011001 10110011001 01110011001 01110011001 11110011001 00001011001 10001011001 01001011001 11001011001 11001011001 00101011001 10101011001 01101011001 11101011001 11101011001 00011011001 10011011001 01011011001 11011011001 11011011001 00111011001 10111011001 01111011001 11111011001 00000111001 00000111001 10000111001 01000111001 11000111001 00100111001 00100111001 10100111001 01100111001 11100111001 00010111001 00010111001 10010111001 01010111001 11010111001 00110111001 00110111001 10110111001 01110111001 11110111001 00001111001 00001111001 10001111001 01001111001 11001111001 00101111001 00101111001 10101111001 01101111001 11101111001 00011111001 00011111001 10011111001 01011111001 11011111001 11011111001 00111111001 10111111001 01111111001 11111111001 11111111001 00000000101 10000000101 01000000101 11000000101 11000000101 00100000101 10100000101 01100000101 01100000101 11100000101 00010000101 10010000101 01010000101 01010000101 11010000101 00110000101 10110000101 10110000101 01110000101 11110000101 00001000101 10001000101 10001000101 01001000101 11001000101 00101000101 00101000101 10101000101 01101000101 11101000101 00011000101 00011000101 10011000101 01011000101 11011000101 11011000101 00111000101 10111000101 01111000101 01111000101 11111000101 00000100101 10000100101 10000100101 01000100101 11000100101 00100100101 10100100101 10100100101 01100100101 11100100101 00010100101 00010100101 10010100101 01010100101 11010100101 11010100101 00110100101 10110100101 01110100101 01110100101 11110100101 00001100101 10001100101 10001100101 01001100101 11001100101 00101100101 00101100101 10101100101 01101100101 11101100101 11101100101 00011100101 10011100101 01011100101 01011100101 11011100101 00111100101 00111100101 10111100101 01111100101 11111100101 11111100101 00000010101 10000010101 01000010101 01000010101 11000010101 00100010101 10100010101 10100010101 01100010101 11100010101 00010010101 00010010101 10010010101 01010010101 01010010101 11010010101 00110010101 10110010101 10110010101 01110010101 11110010101 00001010101 00001010101 10001010101 01001010101 01001010101 11001010101 00101010101 10101010101 10101010101 01101010101 11101010101 11101010101 00011010101 10011010101 01011010101 01011010101 11011010101 00111010101 00111010101 10111010101 01111010101 11111010101 11111010101 00000110101 10000110101 10000110101 01000110101 11000110101 00100110101 00100110101 10100110101 01100110101 01100110101 11100110101 00010110101 10010110101 10010110101 01010110101 11010110101 11010110101 00110110101 10110110101 10110110101 01110110101 11110110101 00001110101 00001110101 10001110101 01001110101 01001110101 11001110101 00101110101 00101110101 10101110101 01101110101 01101110101 11101110101 00011110101 10011110101 10011110101 01011110101 11011110101 11011110101 00111110101 10111110101 10111110101 01111110101 11111110101 11111110101 00000001101 10000001101 10000001101 01000001101 11000001101 11000001101 00100001101 10100001101 01100001101 01100001101 11100001101 00010001101 00010001101 10010001101 01010001101 01010001101 11010001101 00110001101 00110001101 10110001101 01110001101 01110001101 11110001101 00001001101 00001001101 10001001101 01001001101 01001001101 11001001101 00101001101 00101001101 10101001101 01101001101 01101001101 11101001101 00011001101 00011001101 10011001101 01011001101 01011001101 11011001101 00111001101 00111001101 10111001101 01111001101 01111001101 11111001101 11111001101 00000101101 10000101101 10000101101 01000101101 11000101101 11000101101 00100101101 10100101101 10100101101 01100101101 11100101101 11100101101 00010101101 10010101101 10010101101 01010101101 01010101101 11010101101 00110101101 00110101101 10110101101 01110101101 01110101101 11110101101 00001101101 00001101101 10001101101 10001101101 01001101101 11001101101 11001101101 00101101101 10101101101 10101101101 01101101101 11101101101 11101101101 00011101101 00011101101 10011101101 01011101101 01011101101 11011101101 00111101101 00111101101 10111101101 10111101101 01111101101 11111101101 11111101101 00000011101 10000011101 10000011101 01000011101 01000011101 11000011101 00100011101 00100011101 10100011101 10100011101 01100011101 11100011101 11100011101 00010011101 10010011101 10010011101 01010011101 01010011101 11010011101 00110011101 00110011101 10110011101 10110011101 01110011101 11110011101 11110011101 00001011101 00001011101 10001011101 01001011101 01001011101 11001011101 11001011101 00101011101 10101011101 10101011101 01101011101 01101011101 11101011101 00011011101 00011011101 10011011101 10011011101 01011011101 01011011101 11011011101 00111011101 00111011101 10111011101 10111011101 01111011101 11111011101 11111011101 00000111101 00000111101 10000111101 01000111101 01000111101 11000111101 11000111101 00100111101 00100111101 10100111101 01100111101 01100111101 11100111101 11100111101 00010111101 00010111101 10010111101 01010111101 01010111101 11010111101 11010111101 00110111101 00110111101 10110111101 01110111101 01110111101 11110111101 11110111101 00001111101 00001111101 10001111101 01001111101 01001111101 11001111101 11001111101 00101111101 00101111101 10101111101 10101111101 01101111101 11101111101 11101111101 00011111101 00011111101 10011111101 10011111101 01011111101 01011111101 11011111101 00111111101 00111111101 10111111101 10111111101 01111111101 01111111101 11111111101 11111111101 00000000011 00000000011 10000000011 01000000011 01000000011 11000000011 11000000011 00100000011 00100000011 10100000011 10100000011 01100000011 01100000011 11100000011 11100000011 00010000011 10010000011 10010000011 01010000011 01010000011 11010000011 11010000011 00110000011 00110000011 10110000011 10110000011 01110000011 01110000011 11110000011 11110000011 00001000011 00001000011 10001000011 10001000011 01001000011 01001000011 11001000011 00101000011 00101000011 10101000011 10101000011 01101000011 01101000011 11101000011 11101000011 00011000011 00011000011 10011000011 10011000011 01011000011 01011000011 11011000011 11011000011 00111000011 00111000011 10111000011 10111000011 01111000011 01111000011 11111000011 11111000011 00000100011 00000100011 10000100011 10000100011 01000100011 01000100011 11000100011 11000100011 00100100011 00100100011 10100100011 10100100011 01100100011 01100100011 11100100011 11100100011 00010100011 00010100011 10010100011 10010100011 01010100011 01010100011 11010100011 11010100011 00110100011 00110100011 00110100011 10110100011 10110100011 01110100011 01110100011 11110100011 11110100011 00001100011 00001100011 10001100011 10001100011 01001100011 01001100011 11001100011 11001100011 00101100011 00101100011 10101100011 10101100011 10101100011 01101100011 01101100011 11101100011 11101100011 00011100011 00011100011 10011100011 10011100011 01011100011 01011100011 11011100011 11011100011 11011100011 00111100011 00111100011 10111100011 10111100011 01111100011 01111100011 11111100011 11111100011 00000010011 00000010011 00000010011 10000010011 10000010011 01000010011 01000010011 11000010011 11000010011 00100010011 00100010011 00100010011 10100010011 10100010011 01100010011 01100010011 11100010011 11100010011 00010010011 00010010011 00010010011 10010010011 10010010011 01010010011 01010010011 11010010011 11010010011 11010010011 00110010011 00110010011 10110010011 10110010011 01110010011 01110010011 01110010011 11110010011 11110010011 00001010011 00001010011 10001010011 10001010011 10001010011 01001010011 01001010011 11001010011 11001010011 11001010011 00101010011 00101010011 10101010011 10101010011 01101010011 01101010011 01101010011 11101010011 11101010011 00011010011 00011010011 00011010011 10011010011 10011010011 01011010011 01011010011 01011010011 11011010011 11011010011 00111010011 00111010011 00111010011 10111010011 10111010011 01111010011 01111010011 01111010011 11111010011 11111010011 00000110011 00000110011 00000110011 10000110011 10000110011 01000110011 01000110011 01000110011 11000110011 11000110011 11000110011 00100110011 00100110011 10100110011 10100110011 10100110011 01100110011 01100110011 11100110011 11100110011 11100110011 00010110011 00010110011 00010110011 10010110011 10010110011 01010110011 01010110011 01010110011 11010110011 11010110011 11010110011 00110110011 00110110011 00110110011 10110110011 10110110011 01110110011 01110110011 01110110011 11110110011 11110110011 11110110011 00001110011 00001110011 00001110011 10001110011 10001110011 10001110011 01001110011 01001110011 11001110011 11001110011 11001110011 00101110011 00101110011 00101110011 10101110011 10101110011 10101110011 01101110011 01101110011 01101110011 11101110011 11101110011 11101110011 00011110011 00011110011 00011110011 10011110011 10011110011 10011110011 01011110011 01011110011 01011110011 11011110011 11011110011 11011110011 00111110011 00111110011 00111110011 10111110011 10111110011 10111110011 01111110011 01111110011 01111110011 11111110011 11111110011 11111110011 00000001011 00000001011 00000001011 10000001011 10000001011 10000001011 01000001011 01000001011 01000001011 11000001011 11000001011 11000001011 11000001011 00100001011 00100001011 00100001011 10100001011 10100001011 10100001011 01100001011 01100001011 01100001011 11100001011 11100001011 11100001011 11100001011 00010001011 00010001011 00010001011 10010001011 10010001011 10010001011 10010001011 01010001011 01010001011 01010001011 11010001011 11010001011 11010001011 00110001011 00110001011 00110001011 00110001011 10110001011 10110001011 10110001011 01110001011 01110001011 01110001011 01110001011 11110001011 11110001011 11110001011 11110001011 00001001011 00001001011 00001001011 10001001011 10001001011 10001001011 10001001011 01001001011 01001001011 01001001011 01001001011 11001001011 11001001011 11001001011 00101001011 00101001011 00101001011 00101001011 10101001011 10101001011 10101001011 10101001011 01101001011 01101001011 01101001011 01101001011 11101001011 11101001011 11101001011 11101001011 00011001011 00011001011 00011001011 00011001011 10011001011 10011001011 10011001011 10011001011 01011001011 01011001011 01011001011 01011001011 11011001011 11011001011 11011001011 11011001011 00111001011 00111001011 00111001011 00111001011 00111001011 10111001011 10111001011 10111001011 10111001011 01111001011 01111001011 01111001011 01111001011 11111001011 11111001011 11111001011 11111001011 11111001011 00000101011 00000101011 00000101011 00000101011 10000101011 10000101011 10000101011 10000101011 10000101011 01000101011 01000101011 01000101011 01000101011 11000101011 11000101011 11000101011 11000101011 11000101011 00100101011 00100101011 00100101011 00100101011 00100101011 10100101011 10100101011 10100101011 10100101011 10100101011 01100101011 01100101011 01100101011 01100101011 01100101011 11100101011 11100101011 11100101011 11100101011 11100101011 00010101011 00010101011 00010101011 00010101011 00010101011 00010101011 10010101011 10010101011 10010101011 10010101011 10010101011 01010101011 01010101011 01010101011 01010101011 01010101011 01010101011 11010101011 11010101011 11010101011 11010101011 11010101011 11010101011 00110101011 00110101011 00110101011 00110101011 00110101011 00110101011 10110101011 10110101011 10110101011 10110101011 10110101011 10110101011 01110101011 01110101011 01110101011 01110101011 01110101011 01110101011 11110101011 11110101011 11110101011 11110101011 11110101011 11110101011 11110101011 00001101011 00001101011 00001101011 00001101011 00001101011 00001101011 00001101011 10001101011 10001101011 10001101011 10001101011 10001101011 10001101011 10001101011 01001101011 01001101011 01001101011 01001101011 01001101011 01001101011 01001101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 00111101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 11011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 01011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 10011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 00011101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 11101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 01101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 10101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 00101101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 11001101011 01001101011 01001101011 01001101011 01001101011 01001101011 01001101011 01001101011 10001101011 10001101011 10001101011 10001101011 10001101011 10001101011 10001101011 00001101011 00001101011 00001101011 00001101011 00001101011 00001101011 00001101011 11110101011 11110101011 11110101011 11110101011 11110101011 11110101011 01110101011 01110101011 01110101011 01110101011 01110101011 01110101011 10110101011 10110101011 10110101011 10110101011 10110101011 10110101011 00110101011 00110101011 00110101011 00110101011 00110101011 00110101011 11010101011 11010101011 11010101011 11010101011 11010101011 11010101011 01010101011 01010101011 01010101011 01010101011 01010101011 10010101011 10010101011 10010101011 10010101011 10010101011 00010101011 00010101011 00010101011 00010101011 00010101011 11100101011 11100101011 11100101011 11100101011 11100101011 01100101011 01100101011 01100101011 01100101011 01100101011 10100101011 10100101011 10100101011 10100101011 10100101011 00100101011 00100101011 00100101011 00100101011 00100101011 11000101011 11000101011 11000101011 11000101011 01000101011 01000101011 01000101011 01000101011 01000101011 10000101011 10000101011 10000101011 10000101011 00000101011 00000101011 00000101011 00000101011 11111001011 11111001011 11111001011 11111001011 11111001011 01111001011 01111001011 01111001011 01111001011 10111001011 10111001011 10111001011 10111001011 00111001011 00111001011 00111001011 00111001011 11011001011 11011001011 11011001011 11011001011 01011001011 01011001011 01011001011 01011001011 10011001011 10011001011 10011001011 00011001011 00011001011 00011001011 00011001011 11101001011 11101001011 11101001011 11101001011 01101001011 01101001011 01101001011 01101001011 10101001011 10101001011 10101001011 00101001011 00101001011 00101001011 00101001011 11001001011 11001001011 11001001011 01001001011 01001001011 01001001011 01001001011 10001001011 10001001011 10001001011 00001001011 00001001011 00001001011 00001001011 11110001011 11110001011 11110001011 01110001011 01110001011 01110001011 10110001011 10110001011 10110001011 10110001011 00110001011 00110001011 00110001011 11010001011 11010001011 11010001011 01010001011 01010001011 01010001011 10010001011 10010001011 10010001011 10010001011 00010001011 00010001011 00010001011 11100001011 11100001011 11100001011 01100001011 01100001011 01100001011 10100001011 10100001011 10100001011 00100001011 00100001011 00100001011 11000001011 11000001011 11000001011 01000001011 01000001011 01000001011 10000001011 10000001011 10000001011 00000001011 00000001011 00000001011 11111110011 11111110011 11111110011 01111110011 01111110011 10111110011 10111110011 10111110011 00111110011 00111110011 00111110011 11011110011 11011110011 11011110011 01011110011 01011110011 01011110011 10011110011 10011110011 00011110011 00011110011 00011110011 11101110011 11101110011 11101110011 01101110011 01101110011 10101110011 10101110011 10101110011 00101110011 00101110011 00101110011 11001110011 11001110011 01001110011 01001110011 01001110011 10001110011 10001110011 00001110011 00001110011 00001110011 11110110011 11110110011 11110110011 01110110011 01110110011 10110110011 10110110011 10110110011 00110110011 00110110011 11010110011 11010110011 11010110011 01010110011 01010110011 10010110011 10010110011 10010110011 00010110011 00010110011 11100110011 11100110011 01100110011 01100110011 01100110011 10100110011 10100110011 00100110011 00100110011 00100110011 11000110011 11000110011 01000110011 01000110011 10000110011 10000110011 10000110011 00000110011 00000110011 11111010011 11111010011 01111010011 01111010011 01111010011 10111010011 10111010011 00111010011 00111010011 11011010011 11011010011 01011010011 01011010011 01011010011 10011010011 10011010011 00011010011 00011010011 11101010011 11101010011 01101010011 01101010011 01101010011 10101010011 10101010011 00101010011 00101010011 11001010011 11001010011 01001010011 01001010011 10001010011 10001010011 00001010011 00001010011 00001010011 11110010011 11110010011 01110010011 01110010011 10110010011 10110010011 00110010011 00110010011 11010010011 11010010011 01010010011 01010010011 10010010011 10010010011 00010010011 00010010011 11100010011 11100010011 01100010011 01100010011 10100010011 10100010011 00100010011 00100010011 11000010011 11000010011 01000010011 01000010011 10000010011 10000010011 00000010011 00000010011 11111100011 11111100011 01111100011 01111100011 10111100011 10111100011 00111100011 00111100011 11011100011 11011100011 01011100011 01011100011 10011100011 10011100011 00011100011 00011100011 11101100011 11101100011 01101100011 01101100011 10101100011 10101100011 00101100011 00101100011 11001100011 11001100011 01001100011 01001100011 10001100011 00001100011 00001100011 11110100011 11110100011 01110100011 01110100011 10110100011 10110100011 00110100011 00110100011 11010100011 11010100011 01010100011 10010100011 10010100011 00010100011 00010100011 11100100011 11100100011 01100100011 01100100011 10100100011 00100100011 00100100011 11000100011 11000100011 01000100011 01000100011 10000100011 10000100011 00000100011 11111000011 11111000011 01111000011 01111000011 10111000011 10111000011 00111000011 11011000011 11011000011 01011000011 01011000011 10011000011 00011000011 00011000011 11101000011 11101000011 01101000011 01101000011 10101000011 00101000011 00101000011 11001000011 11001000011 01001000011 10001000011 10001000011 00001000011 00001000011 11110000011 01110000011 01110000011 10110000011 10110000011 00110000011 11010000011 11010000011 01010000011 01010000011 10010000011 00010000011 00010000011 11100000011 11100000011 01100000011 10100000011 10100000011 00100000011 00100000011 11000000011 01000000011 01000000011 10000000011 00000000011 00000000011 11111111101 11111111101 01111111101 10111111101 10111111101 00111111101 11011111101 11011111101 01011111101 10011111101 10011111101 00011111101 00011111101 11101111101 01101111101 01101111101 10101111101 00101111101 00101111101 11001111101 01001111101 01001111101 10001111101 00001111101 00001111101 11110111101 11110111101 01110111101 10110111101 10110111101 00110111101 11010111101 11010111101 01010111101 10010111101 10010111101 00010111101 11100111101 11100111101 01100111101 10100111101 10100111101 00100111101 11000111101 11000111101 01000111101 10000111101 10000111101 00000111101 11111011101 11111011101 01111011101 10111011101 00111011101 00111011101 11011011101 01011011101 01011011101 10011011101 00011011101 00011011101 11101011101 01101011101 01101011101 10101011101 00101011101 00101011101 11001011101 01001011101 10001011101 10001011101 00001011101 11110011101 11110011101 01110011101 10110011101 00110011101 00110011101 11010011101 01010011101 01010011101 10010011101 00010011101 00010011101 11100011101 01100011101 10100011101 10100011101 00100011101 11000011101 01000011101 01000011101 10000011101 00000011101 00000011101 11111101101 01111101101 10111101101 10111101101 00111101101 11011101101 01011101101 01011101101 10011101101 00011101101 11101101101 11101101101 01101101101 10101101101 10101101101 00101101101 11001101101 01001101101 01001101101 10001101101 00001101101 11110101101 11110101101 01110101101 10110101101 00110101101 00110101101 11010101101 01010101101 10010101101 00010101101 00010101101 11100101101 01100101101 10100101101 10100101101 00100101101 11000101101 01000101101 01000101101 10000101101 00000101101 11111001101 01111001101 01111001101 10111001101 00111001101 11011001101 11011001101 01011001101 10011001101 00011001101 11101001101 11101001101 01101001101 10101001101 00101001101 11001001101 11001001101 01001001101 10001001101 00001001101 11110001101 11110001101 01110001101 10110001101 00110001101 11010001101 11010001101 01010001101 10010001101 00010001101 11100001101 11100001101 01100001101 10100001101 00100001101 11000001101 11000001101 01000001101 10000001101 00000001101 11111110101 01111110101 01111110101 10111110101 00111110101 11011110101 01011110101 01011110101 10011110101 00011110101 11101110101 01101110101 10101110101 10101110101 00101110101 11001110101 01001110101 10001110101 00001110101 00001110101 11110110101 01110110101 10110110101 00110110101 11010110101 01010110101 01010110101 10010110101 00010110101 11100110101 01100110101 10100110101 00100110101 00100110101 11000110101 01000110101 10000110101 00000110101 11111010101 01111010101 01111010101 10111010101 00111010101 11011010101 01011010101 10011010101 00011010101 00011010101 11101010101 01101010101 10101010101 00101010101 11001010101 01001010101 10001010101 10001010101 00001010101 11110010101 01110010101 10110010101 00110010101 11010010101 01010010101 10010010101 10010010101 00010010101 11100010101 01100010101 10100010101 00100010101 11000010101 01000010101 10000010101 00000010101 00000010101 11111100101 01111100101 10111100101 00111100101 11011100101 01011100101 10011100101 00011100101 11101100101 01101100101 01101100101 10101100101 00101100101 11001100101 01001100101 10001100101 00001100101 11110100101 01110100101 10110100101 00110100101 11010100101 01010100101 01010100101 10010100101 00010100101 11100100101 01100100101 10100100101 00100100101 11000100101 01000100101 10000100101 00000100101 11111000101 01111000101 10111000101 00111000101 11011000101 11011000101 01011000101 10011000101 00011000101 11101000101 01101000101 10101000101 00101000101 11001000101 01001000101 10001000101 00001000101 11110000101 01110000101 10110000101 00110000101 11010000101 01010000101 10010000101 00010000101 11100000101 01100000101 10100000101 00100000101 11000000101 01000000101 10000000101 00000000101 00000000101 11111111001 01111111001 10111111001 00111111001 11011111001 01011111001 10011111001 00011111001 11101111001 01101111001 10101111001 00101111001 11001111001 01001111001 10001111001 00001111001 11110111001 01110111001 10110111001 00110111001 11010111001 01010111001 10010111001 00010111001 11100111001 01100111001 10100111001 00100111001 11000111001 01000111001 10000111001 00000111001 11111011001 01111011001 00111011001 11011011001 01011011001 10011011001 00011011001 11101011001 01101011001 10101011001 00101011001 11001011001 01001011001 10001011001 00001011001 11110011001 01110011001 10110011001 00110011001 11010011001 01010011001 10010011001 00010011001 11100011001 01100011001 10100011001 00100011001 11000011001 01000011001 10000011001 11111101001 01111101001 10111101001 00111101001 11011101001 01011101001 10011101001 00011101001 11101101001 01101101001 10101101001 00101101001 11001101001 01001101001 10001101001 00001101001 01110101001 10110101001 00110101001 11010101001 01010101001 10010101001 00010101001 11100101001 01100101001 10100101001 00100101001 11000101001 01000101001 00000101001 11111001001 01111001001 10111001001 00111001001 11011001001 01011001001 10011001001 00011001001 11101001001 01101001001 00101001001 11001001001 01001001001 10001001001 00001001001 11110001001 01110001001 10110001001 00110001001 11010001001 10010001001 00010001001 11100001001 01100001001 10100001001 00100001001 11000001001 01000001001 00000001001 11111110001 01111110001 10111110001 00111110001 11011110001 01011110001 10011110001 00011110001 01101110001 10101110001 00101110001 11001110001 01001110001 10001110001 00001110001 01110110001 10110110001 00110110001 11010110001 01010110001 10010110001 00010110001 01100110001 10100110001 00100110001 11000110001 01000110001 10000110001 00000110001 01111010001 10111010001 00111010001 11011010001 01011010001 10011010001 11101010001 01101010001 10101010001 00101010001 11001010001 01001010001 00001010001 11110010001 01110010001 10110010001 00110010001 11010010001 10010010001 00010010001 11100010001 01100010001 10100010001 00100010001 01000010001 10000010001 00000010001 11111100001 01111100001 00111100001 11011100001 01011100001 10011100001 00011100001 01101100001 10101100001 00101100001 11001100001 01001100001 10001100001 11110100001 01110100001 10110100001 00110100001 01010100001 10010100001 00010100001 11100100001 01100100001 00100100001 11000100001 01000100001 10000100001 00000100001 01111000001 10111000001 00111000001 11011000001 01011000001 00011000001 11101000001 01101000001 10101000001 11001000001 01001000001 10001000001 00001000001 01110000001 10110000001 00110000001 11010000001 01010000001 00010000001 11100000001 01100000001 10100000001 11000000001 01000000001 10000000001 00000000001 01111111110 10111111110 00111111110 11011111110 10011111110 00011111110 11101111110 01101111110 00101111110 11001111110 01001111110 10001111110 11110111110 01110111110 10110111110 00110111110 01010111110 10010111110 00010111110 01100111110 10100111110 00100111110 11000111110 10000111110 00000111110 11111011110 01111011110 00111011110 11011011110 01011011110 00011011110 11101011110 01101011110 10101011110 11001011110 01001011110 10001011110 11110011110 01110011110 10110011110 00110011110 01010011110 10010011110 00010011110 01100011110 10100011110 00100011110 01000011110 10000011110 00000011110 11111101110 10111101110 00111101110 11011101110 10011101110 00011101110 11101101110 10101101110 00101101110 11001101110 10001101110 00001101110 11110101110 10110101110 00110101110 11010101110 10010101110 00010101110 11100101110 10100101110 00100101110 11000101110 01000101110 00000101110 11111001110 01111001110 00111001110 11011001110 10011001110 00011001110 11101001110 10101001110 00101001110 11001001110 10001001110 00001001110 11110001110 10110001110 00110001110 11010001110 10010001110 00010001110 11100001110 10100001110 00100001110 11000001110 10000001110 00000001110 01111110110 10111110110 00111110110 01011110110 10011110110 00011110110 01101110110 10101110110 00101110110 01001110110 10001110110 11110110110 01110110110 10110110110 11010110110 01010110110 10010110110 11100110110 01100110110 00100110110 11000110110 01000110110 00000110110 11111010110 10111010110 00111010110 11011010110 10011010110 00011010110 01101010110 10101010110 00101010110 01001010110 10001010110 11110010110 01110010110 10110010110 11010010110 01010010110 00010010110 11100010110 01100010110 00100010110 11000010110 10000010110 00000010110 11111100110 10111100110 00111100110 01011100110 10011100110 11101100110 01101100110 10101100110 11001100110 01001100110 00001100110 11110100110 10110100110 00110100110 11010100110 10010100110 00010100110 01100100110 10100100110 11000100110 01000100110 10000100110 11111000110 01111000110 00111000110 11011000110 10011000110 00011000110 01101000110 10101000110 00101000110 01001000110 10001000110 11110000110 01110000110 00110000110 11010000110 10010000110 00010000110 01100000110 10100000110 11000000110 01000000110 10000000110 11111111010 01111111010 00111111010 11011111010 10011111010 00011111010 01101111010 10101111010 11001111010 01001111010 00001111010 11110111010 10110111010 00110111010 01010111010 10010111010 11100111010 01100111010 00100111010 11000111010 10000111010 00000111010 01111011010 10111011010 11011011010 01011011010 00011011010 11101011010 10101011010 00101011010 01001011010 10001011010 11110011010 01110011010 00110011010 11010011010 10010011010 00010011010 01100011010 10100011010 11000011010 01000011010 00000011010 11111101010 10111101010 00111101010 01011101010 10011101010 11101101010 01101101010 00101101010 11001101010 10001101010 00001101010 01110101010 00110101010 11010101010 10010101010 00010101010 01100101010 10100101010 11000101010 01000101010 00000101010 11111001010 10111001010 00111001010 01011001010 00011001010 11101001010 10101001010 00101001010 01001001010 10001001010 11110001010 01110001010 00110001010 01010001010 10010001010 11100001010 01100001010 00100001010 11000001010 10000001010 11111110010 01111110010 00111110010 11011110010 10011110010 00011110010 01101110010 00101110010 11001110010 10001110010 00001110010 01110110010 10110110010 11010110010 10010110010 00010110010 01100110010 10100110010 11000110010 10000110010 00000110010 01111010010 10111010010 11011010010 10011010010 00011010010 01101010010 10101010010 11001010010 10001010010 00001010010 01110010010 10110010010 11010010010 10010010010 00010010010 01100010010 10100010010 11000010010 10000010010 00000010010 01111100010 10111100010 11011100010 10011100010 00011100010 01101100010 00101100010 11001100010 10001100010 00001100010 01110100010 00110100010 11010100010 10010100010 11100100010 01100100010 00100100010 01000100010 10000100010 11111000010 01111000010 00111000010 01011000010 10011000010 11101000010 10101000010 00101000010 01001000010 00001000010 11110000010 10110000010 11010000010 01010000010 00010000010 01100000010 10100000010 11000000010 10000000010 00000000010 01111111100 00111111100 11011111100 10011111100 11101111100 01101111100 00101111100 01001111100 10001111100 11110111100 10110111100 00110111100 01010111100 00010111100 11100111100 10100111100 11000111100 01000111100 00000111100 01111011100 10111011100 11011011100 10011011100 00011011100 01101011100 00101011100 01001011100 10001011100 11110011100 10110011100 00110011100 01010011100 00010011100 11100011100 10100011100 11000011100 10000011100 00000011100 01111101100 00111101100 11011101100 10011101100 11101101100 10101101100 00101101100 01001101100 00001101100 11110101100 10110101100 11010101100 10010101100 00010101100 01100101100 00100101100 11000101100 10000101100 11111001100 10111001100 00111001100 01011001100 00011001100 01101001100 10101001100 11001001100 10001001100 11110001100 01110001100 00110001100 01010001100 00010001100 11100001100 10100001100 11000001100 10000001100 00000001100 01111110100 00111110100 01011110100 10011110100 11101110100 10101110100 11001110100 01001110100 00001110100 01110110100 00110110100 11010110100 10010110100 11100110100 10100110100 11000110100 01000110100 00000110100 01111010100 00111010100 11011010100 10011010100 11101010100 10101010100 11001010100 01001010100 00001010100 01110010100 00110010100 11010010100 10010010100 11100010100 10100010100 11000010100 01000010100 00000010100 01111100100 00111100100 01011100100 10011100100 11101100100 10101100100 11001100100 10001100100 00001100100 01110100100 00110100100 01010100100 00010100100 11100100100 10100100100 11000100100 10000100100 11111000100 10111000100 00111000100 01011000100 00011000100 01101000100 00101000100 11001000100 10001000100 11110000100 10110000100 11010000100 10010000100 00010000100 01100000100 00100000100 01000000100 00000000100 01111111000 10111111000 11011111000 10011111000 11101111000 10101111000 11001111000 10001111000 00001111000 01110111000 00110111000 01010111000 00010111000 01100111000 00100111000 11000111000 10000111000 11111011000 10111011000 11011011000 10011011000 11101011000 01101011000 00101011000 01001011000 00001011000 01110011000 00110011000 01010011000 00010011000 11100011000 10100011000 11000011000 10000011000 11111101000 10111101000 11011101000 10011101000 00011101000 01101101000 00101101000 01001101000 00001101000 01110101000 00110101000 01010101000 00010101000 11100101000 10100101000 11000101000 10000101000 11111001000 10111001000 11011001000 10011001000 11101001000 10101001000 00101001000 01001001000 00001001000 01110001000 00110001000 01010001000 00010001000 01100001000 00100001000 01000001000 00000001000 01111110000 10111110000 11011110000 10011110000 11101110000 10101110000 11001110000 10001110000 11110110000 10110110000 11010110000 10010110000 11100110000 10100110000 11000110000 10000110000 00000110000 01111010000 00111010000 01011010000 00011010000 01101010000 00101010000 01001010000 00001010000 01110010000 00110010000 01010010000 00010010000 01100010000 00100010000 01000010000 00000010000 01111100000 00111100000 01011100000 00011100000 11101100000 10101100000 11001100000 10001100000 11110100000 10110100000 11010100000 10010100000 11100100000 10100100000 11000100000 10000100000 11111000000 10111000000 11011000000 10011000000 11101000000 10101000000 11001000000 10001000000 11110000000 10110000000 11010000000 10010000000 11100000000 10100000000 11000000000 10000000000"),
    .MODE("DP"),
    .OREGSET_A("RESET"),
    .OREGSET_B("RESET"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE_A("ASYNC"),
    .RESETMODE_B("ASYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    al_82f1a528 (
    .addra(al_a07945e6),
    .addrb({al_bf62f43[11:1],al_a07945e6[0]}),
    .bea(1'b0),
    .beb(1'b0),
    .cea(1'b1),
    .ceb(1'b1),
    .clka(clk),
    .clkb(clk),
    .dia(11'b00000000000),
    .dib(11'b00000000000),
    .ocea(1'b1),
    .oceb(1'b1),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(1'b0),
    .web(1'b0),
    .doa(al_80d2564a),
    .dob(al_8aaaf100));
  AL_DFF_X al_dcfce2f0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(1'b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25fbcbb5));
  AL_DFF_X al_81c3b7c8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_25fbcbb5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(rdy));
  AL_DFF_X al_e2342da (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[8]));
  AL_DFF_X al_f8c23993 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[9]));
  AL_DFF_X al_7f0c0435 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[10]));
  AL_DFF_X al_b354880f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[11]));
  AL_DFF_X al_b3ef0560 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[12]));
  AL_DFF_X al_a0292264 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[13]));
  AL_DFF_X al_ac9b3078 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[14]));
  AL_DFF_X al_fd18d67 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[15]));
  AL_DFF_X al_d6bb0029 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[16]));
  AL_DFF_X al_474f8f4a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[17]));
  AL_DFF_X al_b26d62bf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[0]));
  AL_DFF_X al_ab9dd774 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[18]));
  AL_DFF_X al_88b39ea0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[19]));
  AL_DFF_X al_9db2f7ba (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[20]));
  AL_DFF_X al_4354aafd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[21]));
  AL_DFF_X al_ab055865 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[22]));
  AL_DFF_X al_9f75260d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[23]));
  AL_DFF_X al_aa1e0ec3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[24]));
  AL_DFF_X al_e9f72998 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[25]));
  AL_DFF_X al_3d07ae02 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[26]));
  AL_DFF_X al_4f22adc1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[27]));
  AL_DFF_X al_809f7104 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[1]));
  AL_DFF_X al_16a9ca3a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[28]));
  AL_DFF_X al_c0fff07d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[29]));
  AL_DFF_X al_8fe65937 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[30]));
  AL_DFF_X al_65d1adb3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[31]));
  AL_DFF_X al_c1468025 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[2]));
  AL_DFF_X al_c19d8344 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[3]));
  AL_DFF_X al_ca1eda73 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[4]));
  AL_DFF_X al_fa89b429 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[5]));
  AL_DFF_X al_3462fe16 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[6]));
  AL_DFF_X al_87f5414c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7521c31[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c12045b[7]));
  AL_DFF_X al_795dec5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[8]));
  AL_DFF_X al_e8b27f0a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[9]));
  AL_DFF_X al_34c43e91 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[10]));
  AL_DFF_X al_4034d121 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[11]));
  AL_DFF_X al_7260e525 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[12]));
  AL_DFF_X al_6eb318e4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[0]));
  AL_DFF_X al_10074c95 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[1]));
  AL_DFF_X al_5fb1cf51 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[2]));
  AL_DFF_X al_dc5daab3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[3]));
  AL_DFF_X al_5394044a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[4]));
  AL_DFF_X al_b89d9b42 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[5]));
  AL_DFF_X al_81c5ed9a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[6]));
  AL_DFF_X al_9e15c642 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_e1c1520b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75776e99[7]));
  AL_DFF_X al_c26c9bb1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[8]));
  AL_DFF_X al_7256805c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[9]));
  AL_DFF_X al_3579341e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[10]));
  AL_DFF_X al_b7079f11 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[11]));
  AL_DFF_X al_89cb7fac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[12]));
  AL_DFF_X al_7f48cb2c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[13]));
  AL_DFF_X al_8c60f702 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[14]));
  AL_DFF_X al_2e772330 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[15]));
  AL_DFF_X al_835d154d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[16]));
  AL_DFF_X al_d32f36bb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[17]));
  AL_DFF_X al_de040350 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[0]));
  AL_DFF_X al_46b4672d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[18]));
  AL_DFF_X al_e10b0f3c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[19]));
  AL_DFF_X al_53e9dc14 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[20]));
  AL_DFF_X al_d79ebee3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[21]));
  AL_DFF_X al_f0bb2d9b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[22]));
  AL_DFF_X al_1faffb9a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[23]));
  AL_DFF_X al_ed14148e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[24]));
  AL_DFF_X al_88b7b6db (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[25]));
  AL_DFF_X al_527d2456 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[26]));
  AL_DFF_X al_7e32d61 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[27]));
  AL_DFF_X al_25378cfc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[1]));
  AL_DFF_X al_77d3213b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[28]));
  AL_DFF_X al_a94d40f9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[29]));
  AL_DFF_X al_8ee8ac50 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[30]));
  AL_DFF_X al_5fba7a49 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[31]));
  AL_DFF_X al_dc93576e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[2]));
  AL_DFF_X al_76b20766 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[3]));
  AL_DFF_X al_a8ce422 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[4]));
  AL_DFF_X al_e3895fe2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[5]));
  AL_DFF_X al_2160ccea (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[6]));
  AL_DFF_X al_df8e007c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(fword[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e800bf9[7]));
  AL_DFF_X al_b40a42c0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[8]));
  AL_DFF_X al_56fbb473 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[9]));
  AL_DFF_X al_f912cfa7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[10]));
  AL_DFF_X al_790357b6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[11]));
  AL_DFF_X al_1f745e25 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[12]));
  AL_DFF_X al_fdf3d1b5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[13]));
  AL_DFF_X al_28c56aa6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[14]));
  AL_DFF_X al_fa1f6a4e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[15]));
  AL_DFF_X al_7852efc4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[16]));
  AL_DFF_X al_9a72719d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[17]));
  AL_DFF_X al_31c2c18 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[0]));
  AL_DFF_X al_7eeaf50d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[18]));
  AL_DFF_X al_3b36aef9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[19]));
  AL_DFF_X al_26b87d2b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[20]));
  AL_DFF_X al_8a5c27f2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[21]));
  AL_DFF_X al_45e64a4e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[22]));
  AL_DFF_X al_33b37756 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[23]));
  AL_DFF_X al_de0a6607 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[24]));
  AL_DFF_X al_e5e3578e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[25]));
  AL_DFF_X al_a8a8dd4b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[26]));
  AL_DFF_X al_d9ae9d4c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[27]));
  AL_DFF_X al_bed75354 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[1]));
  AL_DFF_X al_9fa6fc7e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[28]));
  AL_DFF_X al_c3aeda92 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[29]));
  AL_DFF_X al_d8454c67 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[30]));
  AL_DFF_X al_7e8984c3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[31]));
  AL_DFF_X al_b2c2a4b7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[2]));
  AL_DFF_X al_99383aba (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[3]));
  AL_DFF_X al_f8178b2c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[4]));
  AL_DFF_X al_be1fc3e5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[5]));
  AL_DFF_X al_c9f8b2f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[6]));
  AL_DFF_X al_5979435b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ac33d53a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2adbf503[7]));
  AL_DFF_X al_efc104d9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[8]));
  AL_DFF_X al_94d694ac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[9]));
  AL_DFF_X al_35f4ffbe (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[10]));
  AL_DFF_X al_38c08d06 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[11]));
  AL_DFF_X al_b4006c49 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[12]));
  AL_DFF_X al_88983c15 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[13]));
  AL_DFF_X al_322c5a5a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[14]));
  AL_DFF_X al_f7f9a105 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[15]));
  AL_DFF_X al_b6c3af5b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[16]));
  AL_DFF_X al_516abd0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[17]));
  AL_DFF_X al_22aeac4e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[0]));
  AL_DFF_X al_2cfb0659 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[18]));
  AL_DFF_X al_7018cf5a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[19]));
  AL_DFF_X al_665b406a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[20]));
  AL_DFF_X al_dd3c6cbd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[21]));
  AL_DFF_X al_88ad635d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[22]));
  AL_DFF_X al_cc28c7fc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[23]));
  AL_DFF_X al_3a1809be (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[24]));
  AL_DFF_X al_f6441446 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[25]));
  AL_DFF_X al_8863e9a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[26]));
  AL_DFF_X al_5e7497d4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[27]));
  AL_DFF_X al_6d6ea447 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[1]));
  AL_DFF_X al_5209be15 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[28]));
  AL_DFF_X al_442ae8f6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[29]));
  AL_DFF_X al_147a8585 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[30]));
  AL_DFF_X al_718633aa (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[31]));
  AL_DFF_X al_1164b4aa (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[2]));
  AL_DFF_X al_ddd1c04b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[3]));
  AL_DFF_X al_bf982701 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[4]));
  AL_DFF_X al_34da7a0f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[5]));
  AL_DFF_X al_b67c3979 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[6]));
  AL_DFF_X al_7d3b3b7c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2adbf503[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1ca72219[7]));
  AL_DFF_X al_67237772 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[8]));
  AL_DFF_X al_5943f200 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[9]));
  AL_DFF_X al_bd8fdd97 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[10]));
  AL_DFF_X al_b9e3c79f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[11]));
  AL_DFF_X al_ac0bcbeb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[12]));
  AL_DFF_X al_13b0591a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[13]));
  AL_DFF_X al_8f28d3a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[14]));
  AL_DFF_X al_7b5d1323 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[15]));
  AL_DFF_X al_5ce47d62 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[16]));
  AL_DFF_X al_db7ed5ae (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[17]));
  AL_DFF_X al_252ea06e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[0]));
  AL_DFF_X al_b7ce14ac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[18]));
  AL_DFF_X al_24230e71 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[19]));
  AL_DFF_X al_957d5748 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[20]));
  AL_DFF_X al_d5572c6e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[21]));
  AL_DFF_X al_157cd271 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[22]));
  AL_DFF_X al_95d30c7f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[23]));
  AL_DFF_X al_fc015cba (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[24]));
  AL_DFF_X al_5f2f12df (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[25]));
  AL_DFF_X al_578df8e9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[26]));
  AL_DFF_X al_605d9003 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[27]));
  AL_DFF_X al_8e33936e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[1]));
  AL_DFF_X al_fe620a1d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[28]));
  AL_DFF_X al_1cc64d73 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[29]));
  AL_DFF_X al_fd757df4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[30]));
  AL_DFF_X al_17f55510 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[31]));
  AL_DFF_X al_2c9f1ebd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[2]));
  AL_DFF_X al_c05bd12f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[3]));
  AL_DFF_X al_7d49ed41 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[4]));
  AL_DFF_X al_6beff56 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[5]));
  AL_DFF_X al_c4f13542 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[6]));
  AL_DFF_X al_86c33c3f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1ca72219[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc74dd1[7]));
  AL_DFF_X al_6f91b8e8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[8]));
  AL_DFF_X al_10ad84aa (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[9]));
  AL_DFF_X al_46410d76 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[10]));
  AL_DFF_X al_93743f2f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[11]));
  AL_DFF_X al_f1db63d4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[0]));
  AL_DFF_X al_fdf401f2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[1]));
  AL_DFF_X al_123f376 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[2]));
  AL_DFF_X al_c051e0c9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[3]));
  AL_DFF_X al_fb384ab2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[4]));
  AL_DFF_X al_141203dd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[5]));
  AL_DFF_X al_51f4caf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[6]));
  AL_DFF_X al_3e10bc68 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_3bc6703c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_50d27df2[7]));
  AL_DFF_X al_6aaae735 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[8]));
  AL_DFF_X al_99a4dbf1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[9]));
  AL_DFF_X al_d82a3ae1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[10]));
  AL_DFF_X al_8254204c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[11]));
  AL_DFF_X al_a2077ece (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[12]));
  AL_DFF_X al_1a7734a8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[13]));
  AL_DFF_X al_233a96c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[14]));
  AL_DFF_X al_7d0868c5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[15]));
  AL_DFF_X al_9a81103f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[16]));
  AL_DFF_X al_6c10bd3c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[17]));
  AL_DFF_X al_b9877cbc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[0]));
  AL_DFF_X al_197f714d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[19]));
  AL_DFF_X al_a908572e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[20]));
  AL_DFF_X al_89a8492 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[21]));
  AL_DFF_X al_85390814 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[22]));
  AL_DFF_X al_e41b1a3a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[23]));
  AL_DFF_X al_31d3fe88 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[24]));
  AL_DFF_X al_e172090b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[25]));
  AL_DFF_X al_d724aa3d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[26]));
  AL_DFF_X al_84c9934c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[27]));
  AL_DFF_X al_d38326ed (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[1]));
  AL_DFF_X al_83e055a4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[28]));
  AL_DFF_X al_3ba0882a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[29]));
  AL_DFF_X al_6e263ab4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[30]));
  AL_DFF_X al_6d3b1c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[31]));
  AL_DFF_X al_c75b9434 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[2]));
  AL_DFF_X al_23f710d6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[3]));
  AL_DFF_X al_1774ae79 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[4]));
  AL_DFF_X al_8086a947 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[5]));
  AL_DFF_X al_50d71bcf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[6]));
  AL_DFF_X al_2965d8d3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc74dd1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_45f60c58[7]));
  AL_DFF_X al_b40e8e05 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[8]));
  AL_DFF_X al_2259e8d1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[9]));
  AL_DFF_X al_5f624aaf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[10]));
  AL_DFF_X al_fd544ba8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[0]));
  AL_DFF_X al_40ebe0d4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[1]));
  AL_DFF_X al_b4cd3408 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[2]));
  AL_DFF_X al_16607eff (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[3]));
  AL_DFF_X al_2e1082f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[4]));
  AL_DFF_X al_806f02ed (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[5]));
  AL_DFF_X al_e97bb64b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[6]));
  AL_DFF_X al_f7f2da08 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_80d2564a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35c5bf4a[7]));
  AL_DFF_X al_e913a317 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[8]));
  AL_DFF_X al_b03a90ff (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[9]));
  AL_DFF_X al_6affaeca (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[10]));
  AL_DFF_X al_60890717 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[11]));
  AL_DFF_X al_bc18c7fd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_50d27df2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[0]));
  AL_DFF_X al_96f1f8a7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[1]));
  AL_DFF_X al_fca51337 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[2]));
  AL_DFF_X al_3957d799 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[3]));
  AL_DFF_X al_755dd614 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[4]));
  AL_DFF_X al_b2433da2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[5]));
  AL_DFF_X al_a11536f6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[6]));
  AL_DFF_X al_91797866 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ef10e9eb[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a07945e6[7]));
  AL_DFF_X al_62640248 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[8]));
  AL_DFF_X al_3ac46452 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[9]));
  AL_DFF_X al_43288d86 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[10]));
  AL_DFF_X al_11932a20 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[11]));
  AL_DFF_X al_5d88f5b2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[12]));
  AL_DFF_X al_7bc6d8aa (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[13]));
  AL_DFF_X al_e235ba43 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[14]));
  AL_DFF_X al_ffa9d9a4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[15]));
  AL_DFF_X al_b5960a71 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[16]));
  AL_DFF_X al_5068432d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[17]));
  AL_DFF_X al_e95fcb14 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[0]));
  AL_DFF_X al_79c45c1a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[19]));
  AL_DFF_X al_4d6db486 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[20]));
  AL_DFF_X al_18688e16 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[21]));
  AL_DFF_X al_484fae1a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[22]));
  AL_DFF_X al_fa83a62b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[23]));
  AL_DFF_X al_fbaceb55 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[24]));
  AL_DFF_X al_569d22f7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[25]));
  AL_DFF_X al_ee584424 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[26]));
  AL_DFF_X al_cd1dc485 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[27]));
  AL_DFF_X al_f488aa32 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[1]));
  AL_DFF_X al_6995a8ac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[28]));
  AL_DFF_X al_412de6e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[29]));
  AL_DFF_X al_552e8945 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[30]));
  AL_DFF_X al_3678cb57 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[31]));
  AL_DFF_X al_a079e3e9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[2]));
  AL_DFF_X al_7d0ad31 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[3]));
  AL_DFF_X al_430c2c91 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[4]));
  AL_DFF_X al_7d86140d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[5]));
  AL_DFF_X al_74e57733 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[6]));
  AL_DFF_X al_bb220e36 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_45f60c58[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf05573[7]));
  AL_DFF_X al_a5f6491e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[8]));
  AL_DFF_X al_4402b56f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[9]));
  AL_DFF_X al_95c0e8ec (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[10]));
  AL_DFF_X al_8a88eb8c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[11]));
  AL_DFF_X al_25e9fff5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[1]));
  AL_DFF_X al_4376c392 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[2]));
  AL_DFF_X al_549078f7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[3]));
  AL_DFF_X al_aa29b77f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[4]));
  AL_DFF_X al_f61e0c79 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[5]));
  AL_DFF_X al_cd459a96 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[6]));
  AL_DFF_X al_9f40c8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_1db9833e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf62f43[7]));
  AL_DFF_X al_f463089f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[8]));
  AL_DFF_X al_6e0c2818 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[9]));
  AL_DFF_X al_7b397e76 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[10]));
  AL_DFF_X al_895e278b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[11]));
  AL_DFF_X al_84ce4441 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[0]));
  AL_DFF_X al_754f7138 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[1]));
  AL_DFF_X al_81333aeb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[2]));
  AL_DFF_X al_9da07d15 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[3]));
  AL_DFF_X al_e8bee181 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[4]));
  AL_DFF_X al_32045acf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[5]));
  AL_DFF_X al_2d1a68c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[6]));
  AL_DFF_X al_1f408e76 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_a07945e6[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aeba03f9[7]));
  AL_DFF_X al_b9f263b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[8]));
  AL_DFF_X al_ef247d1d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[9]));
  AL_DFF_X al_88cef0c5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[10]));
  AL_DFF_X al_38d68827 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[11]));
  AL_DFF_X al_cb3d60b7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[12]));
  AL_DFF_X al_5a147783 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[13]));
  AL_DFF_X al_823353cb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[14]));
  AL_DFF_X al_ce19b6f8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[15]));
  AL_DFF_X al_bad3147f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[16]));
  AL_DFF_X al_ec0bf094 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[17]));
  AL_DFF_X al_87c44ef5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[0]));
  AL_DFF_X al_74272628 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[19]));
  AL_DFF_X al_54dd845a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[20]));
  AL_DFF_X al_6157745c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[21]));
  AL_DFF_X al_1f7bf6af (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[22]));
  AL_DFF_X al_72678665 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[23]));
  AL_DFF_X al_25fc5773 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[24]));
  AL_DFF_X al_216dcd8b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[25]));
  AL_DFF_X al_a9581d71 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[26]));
  AL_DFF_X al_4fd21f4c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[27]));
  AL_DFF_X al_67fe22ba (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[1]));
  AL_DFF_X al_b3fe40f4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[28]));
  AL_DFF_X al_22d1016d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[29]));
  AL_DFF_X al_12edf336 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[30]));
  AL_DFF_X al_b329657a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[31]));
  AL_DFF_X al_e625d767 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[2]));
  AL_DFF_X al_6d1e9f4b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[3]));
  AL_DFF_X al_67d9a12d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[4]));
  AL_DFF_X al_f0e27fb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[5]));
  AL_DFF_X al_5bb451a6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[6]));
  AL_DFF_X al_4b1214b2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf05573[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b84f9223[7]));
  AL_DFF_X al_172e702a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[8]));
  AL_DFF_X al_222268e1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[9]));
  AL_DFF_X al_d547d22d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[10]));
  AL_DFF_X al_a3bae4a6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[11]));
  AL_DFF_X al_44a87bd3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[1]));
  AL_DFF_X al_5db6e7a6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[2]));
  AL_DFF_X al_ce317ef3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[3]));
  AL_DFF_X al_abba78ac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[4]));
  AL_DFF_X al_c6d88610 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[5]));
  AL_DFF_X al_d0603f29 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[6]));
  AL_DFF_X al_f8828ab4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bf62f43[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c65e87[7]));
  AL_DFF_X al_4fc9cae5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[8]));
  AL_DFF_X al_7a12e980 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[9]));
  AL_DFF_X al_7669782b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[10]));
  AL_DFF_X al_4ff3c2ce (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[11]));
  AL_DFF_X al_ac4d7424 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[0]));
  AL_DFF_X al_55c36923 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[1]));
  AL_DFF_X al_193fbe53 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[2]));
  AL_DFF_X al_690bf002 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[3]));
  AL_DFF_X al_85cb4108 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[4]));
  AL_DFF_X al_7146fac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[5]));
  AL_DFF_X al_20c9901f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[6]));
  AL_DFF_X al_43bfe00a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_aeba03f9[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9644e37b[7]));
  AL_DFF_X al_ed1b7004 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[8]));
  AL_DFF_X al_63c28c0e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[9]));
  AL_DFF_X al_8534e5ed (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[10]));
  AL_DFF_X al_e6f668b9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[11]));
  AL_DFF_X al_7fddc7e8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[12]));
  AL_DFF_X al_3e6c67ae (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[13]));
  AL_DFF_X al_e5975af6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[14]));
  AL_DFF_X al_634bfbd2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[15]));
  AL_DFF_X al_ef48f93d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[16]));
  AL_DFF_X al_a0fa41ba (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[17]));
  AL_DFF_X al_66c9a2d5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[0]));
  AL_DFF_X al_b8e08420 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[19]));
  AL_DFF_X al_7beded76 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[20]));
  AL_DFF_X al_999d182f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[21]));
  AL_DFF_X al_91f18bd5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[22]));
  AL_DFF_X al_43e8b10f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[23]));
  AL_DFF_X al_b870df5c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[24]));
  AL_DFF_X al_28492c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[25]));
  AL_DFF_X al_d5d357e2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[26]));
  AL_DFF_X al_f6c31888 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[27]));
  AL_DFF_X al_6e1958fc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[1]));
  AL_DFF_X al_949bcee3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[28]));
  AL_DFF_X al_1e3f5585 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[29]));
  AL_DFF_X al_8f292899 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[30]));
  AL_DFF_X al_559468df (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[31]));
  AL_DFF_X al_effe3088 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[2]));
  AL_DFF_X al_3a5ab10a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[3]));
  AL_DFF_X al_d3492ef6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[4]));
  AL_DFF_X al_622d1db4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[5]));
  AL_DFF_X al_819c9fac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[6]));
  AL_DFF_X al_e9484e4c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b84f9223[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fd1686[7]));
  AL_DFF_X al_d753fd8a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[8]));
  AL_DFF_X al_5838e2a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[9]));
  AL_DFF_X al_65e6ae15 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[10]));
  AL_DFF_X al_37cf9796 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[11]));
  AL_DFF_X al_fef96879 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[1]));
  AL_DFF_X al_6ed237a5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[2]));
  AL_DFF_X al_19c523b2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[3]));
  AL_DFF_X al_6d931c57 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[4]));
  AL_DFF_X al_7874f440 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[5]));
  AL_DFF_X al_e20d8638 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[6]));
  AL_DFF_X al_90c645d6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_2c65e87[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff8d588f[7]));
  AL_DFF_X al_4bd759f7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[8]));
  AL_DFF_X al_e796952d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[9]));
  AL_DFF_X al_f1b26430 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[10]));
  AL_DFF_X al_f9d83a34 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[11]));
  AL_DFF_X al_114d8c6b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[0]));
  AL_DFF_X al_3be727b6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[1]));
  AL_DFF_X al_d1f4536b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[2]));
  AL_DFF_X al_e9a3754d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[3]));
  AL_DFF_X al_d4d3d7b4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[4]));
  AL_DFF_X al_941a71ae (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[5]));
  AL_DFF_X al_af6015e2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[6]));
  AL_DFF_X al_9da12de8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_9644e37b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0376e91[7]));
  AL_DFF_X al_596b0fc4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[8]));
  AL_DFF_X al_5cfa2c1e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[9]));
  AL_DFF_X al_c56c02f8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[10]));
  AL_DFF_X al_16ad90bc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[0]));
  AL_DFF_X al_e1044ec0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[1]));
  AL_DFF_X al_16da6de4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[2]));
  AL_DFF_X al_e819e904 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[3]));
  AL_DFF_X al_4990808d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[4]));
  AL_DFF_X al_d51e17ed (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[5]));
  AL_DFF_X al_b67f884b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[6]));
  AL_DFF_X al_ff3308ea (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_35c5bf4a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b33e7450[7]));
  AL_DFF_X al_6f646297 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[8]));
  AL_DFF_X al_e9f5eab5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[9]));
  AL_DFF_X al_73eb83df (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[10]));
  AL_DFF_X al_2f1827e9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[11]));
  AL_DFF_X al_1f4569df (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[12]));
  AL_DFF_X al_663c9601 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[13]));
  AL_DFF_X al_6d500715 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[14]));
  AL_DFF_X al_a1505949 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[15]));
  AL_DFF_X al_2c6e7404 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[16]));
  AL_DFF_X al_268928b1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[17]));
  AL_DFF_X al_bb8e61f6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[0]));
  AL_DFF_X al_73683ddd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[19]));
  AL_DFF_X al_dbfe227c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[20]));
  AL_DFF_X al_5542e6f4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[21]));
  AL_DFF_X al_a7e1139b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[22]));
  AL_DFF_X al_1409141a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[23]));
  AL_DFF_X al_66ab83d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[24]));
  AL_DFF_X al_53e7291c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[25]));
  AL_DFF_X al_cdcc863a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[26]));
  AL_DFF_X al_ded83a89 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[27]));
  AL_DFF_X al_cac62b2f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[1]));
  AL_DFF_X al_4f4242dc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[28]));
  AL_DFF_X al_e918d966 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[29]));
  AL_DFF_X al_a50abdd1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[30]));
  AL_DFF_X al_ca73761c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[31]));
  AL_DFF_X al_640d9f02 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[2]));
  AL_DFF_X al_57fa46a5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[3]));
  AL_DFF_X al_3e8f5316 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[4]));
  AL_DFF_X al_7fa0bf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[5]));
  AL_DFF_X al_62a03df9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[6]));
  AL_DFF_X al_617dc28a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8fd1686[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fdd6779[7]));
  AL_DFF_X al_e94e1ee5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[8]));
  AL_DFF_X al_41d42908 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[9]));
  AL_DFF_X al_2482afa0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[10]));
  AL_DFF_X al_c191b8f5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[11]));
  AL_DFF_X al_dd12912b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[1]));
  AL_DFF_X al_52a21520 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[2]));
  AL_DFF_X al_484fdc03 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[3]));
  AL_DFF_X al_8cc9e864 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[4]));
  AL_DFF_X al_2f7c5fd5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[5]));
  AL_DFF_X al_e6bf6678 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[6]));
  AL_DFF_X al_4f91ad1f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_ff8d588f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e765e4ce[7]));
  AL_DFF_X al_25497697 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[8]));
  AL_DFF_X al_a6031452 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[9]));
  AL_DFF_X al_a28ca941 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[10]));
  AL_DFF_X al_f33fc8f6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[11]));
  AL_DFF_X al_c07f6b33 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[12]));
  AL_DFF_X al_c520b2e8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[13]));
  AL_DFF_X al_97360cc1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[14]));
  AL_DFF_X al_687ba53e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[15]));
  AL_DFF_X al_259027fb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[16]));
  AL_DFF_X al_33faba75 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[17]));
  AL_DFF_X al_bf6fc322 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[0]));
  AL_DFF_X al_c4008a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b0376e91[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[18]));
  AL_DFF_X al_e84489ed (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[19]));
  AL_DFF_X al_136e443c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[20]));
  AL_DFF_X al_e8ec7a28 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[21]));
  AL_DFF_X al_21e3964 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[22]));
  AL_DFF_X al_a137efc6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[23]));
  AL_DFF_X al_43a6a0c7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[24]));
  AL_DFF_X al_1fa43b18 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[25]));
  AL_DFF_X al_3062ba06 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[26]));
  AL_DFF_X al_67dcc451 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[27]));
  AL_DFF_X al_58ee35ea (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[1]));
  AL_DFF_X al_f82aec5c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[28]));
  AL_DFF_X al_ec3557a6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[29]));
  AL_DFF_X al_12328588 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[30]));
  AL_DFF_X al_3fdac79f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[31]));
  AL_DFF_X al_9f89269f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[2]));
  AL_DFF_X al_fd7fb13b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[3]));
  AL_DFF_X al_64d1e8bd (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[4]));
  AL_DFF_X al_7f86ac5b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[5]));
  AL_DFF_X al_82dfed12 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[6]));
  AL_DFF_X al_3fcdd17c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_4fdd6779[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_411d7869[7]));
  AL_DFF_X al_af1970ee (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[8]));
  AL_DFF_X al_4386b1d1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[9]));
  AL_DFF_X al_39f1326b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[10]));
  AL_DFF_X al_bf5ea2e6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[11]));
  AL_DFF_X al_8474ec3e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[12]));
  AL_DFF_X al_f654e053 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[13]));
  AL_DFF_X al_64a1a276 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[14]));
  AL_DFF_X al_7470868b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[15]));
  AL_DFF_X al_e2f72ab5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[16]));
  AL_DFF_X al_719f4b1c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[17]));
  AL_DFF_X al_ec25c2ce (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[0]));
  AL_DFF_X al_267beac6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[18]));
  AL_DFF_X al_add1732c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[19]));
  AL_DFF_X al_9ff12ce3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[20]));
  AL_DFF_X al_df0357f5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[21]));
  AL_DFF_X al_3dfa252f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[22]));
  AL_DFF_X al_61789b78 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[23]));
  AL_DFF_X al_e6debad6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[24]));
  AL_DFF_X al_824448d9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[25]));
  AL_DFF_X al_72bef55c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[26]));
  AL_DFF_X al_1a00d0bb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[27]));
  AL_DFF_X al_92bcc675 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[1]));
  AL_DFF_X al_c3bafeaf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[28]));
  AL_DFF_X al_80fe0c2a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[29]));
  AL_DFF_X al_1e4e26da (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[30]));
  AL_DFF_X al_ac9f6945 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[31]));
  AL_DFF_X al_eb76298 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[2]));
  AL_DFF_X al_f1e3be7a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[3]));
  AL_DFF_X al_33031e60 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[4]));
  AL_DFF_X al_b4c4dee5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[5]));
  AL_DFF_X al_4b8f3f49 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[6]));
  AL_DFF_X al_d8d633b1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_411d7869[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_347def8c[7]));
  AL_DFF_X al_962d1cf7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[8]));
  AL_DFF_X al_fd50410f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[9]));
  AL_DFF_X al_42e0f270 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[10]));
  AL_DFF_X al_3f1902d2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[11]));
  AL_DFF_X al_b1622de2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[12]));
  AL_DFF_X al_5a5133a3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[13]));
  AL_DFF_X al_b9125c23 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[14]));
  AL_DFF_X al_1c9f534c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[15]));
  AL_DFF_X al_4564e9f9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[16]));
  AL_DFF_X al_1295078 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[17]));
  AL_DFF_X al_209580d8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[0]));
  AL_DFF_X al_3781e35b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[18]));
  AL_DFF_X al_4d62fe79 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[19]));
  AL_DFF_X al_1526c6c7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[20]));
  AL_DFF_X al_49e99c9b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[21]));
  AL_DFF_X al_e18c1919 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[22]));
  AL_DFF_X al_6948eb91 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[23]));
  AL_DFF_X al_95405f63 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[24]));
  AL_DFF_X al_661c41c3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[25]));
  AL_DFF_X al_bc8be88 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[26]));
  AL_DFF_X al_9f722b75 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[27]));
  AL_DFF_X al_6c1e3f36 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[1]));
  AL_DFF_X al_7f6681ac (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[28]));
  AL_DFF_X al_cf5c189e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[29]));
  AL_DFF_X al_312cdcce (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[30]));
  AL_DFF_X al_510b6197 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[31]));
  AL_DFF_X al_6890c3a3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[2]));
  AL_DFF_X al_82fa996c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[3]));
  AL_DFF_X al_17fc00eb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[4]));
  AL_DFF_X al_61d44e82 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[5]));
  AL_DFF_X al_dabba857 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[6]));
  AL_DFF_X al_1806a236 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_347def8c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(phase_out[7]));
  AL_DFF_X al_bbf2313f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[8]));
  AL_DFF_X al_f26ffcf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[9]));
  AL_DFF_X al_540e2433 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[10]));
  AL_DFF_X al_31000d5e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[11]));
  AL_DFF_X al_3b8343fc (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[12]));
  AL_DFF_X al_bd06ff71 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[13]));
  AL_DFF_X al_a9dddd3a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[14]));
  AL_DFF_X al_37d2cf39 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[15]));
  AL_DFF_X al_1032901 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[16]));
  AL_DFF_X al_1f965578 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[17]));
  AL_DFF_X al_f405b828 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[0]));
  AL_DFF_X al_c9dc536d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[18]));
  AL_DFF_X al_c008d929 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[19]));
  AL_DFF_X al_c5f46f5f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[20]));
  AL_DFF_X al_4ad700b0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[21]));
  AL_DFF_X al_47e751e3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[22]));
  AL_DFF_X al_cfdef369 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[23]));
  AL_DFF_X al_44686d66 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[24]));
  AL_DFF_X al_bbcf31b8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[25]));
  AL_DFF_X al_d74a3678 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[26]));
  AL_DFF_X al_4b5ec9a9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[27]));
  AL_DFF_X al_e2c72155 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[1]));
  AL_DFF_X al_e93783b2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[28]));
  AL_DFF_X al_49b895d3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[29]));
  AL_DFF_X al_7ecc318 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[30]));
  AL_DFF_X al_9f9cb2c5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[31]));
  AL_DFF_X al_7dd886c0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[2]));
  AL_DFF_X al_5987efe6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[3]));
  AL_DFF_X al_3daa3114 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[4]));
  AL_DFF_X al_86102fda (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[5]));
  AL_DFF_X al_c9ea4bc7 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[6]));
  AL_DFF_X al_78c44601 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(pword[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2fc0f064[7]));
  AL_DFF_X al_80f3d39a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[8]));
  AL_DFF_X al_601fbdc2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[9]));
  AL_DFF_X al_55318a6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[10]));
  AL_DFF_X al_84118ef1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[11]));
  AL_DFF_X al_4d5bdb82 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[12]));
  AL_DFF_X al_3f441238 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[13]));
  AL_DFF_X al_6752fdd0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_7cb3139[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[0]));
  AL_DFF_X al_7448eb2c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[1]));
  AL_DFF_X al_ddc32b41 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[2]));
  AL_DFF_X al_2df93afe (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[3]));
  AL_DFF_X al_f0c9e6c4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[4]));
  AL_DFF_X al_75b48974 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[5]));
  AL_DFF_X al_f7208ae6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[6]));
  AL_DFF_X al_c0347f07 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6b994b8c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_cos[7]));
  AL_DFF_X al_c49228bf (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[8]));
  AL_DFF_X al_2602aec6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[9]));
  AL_DFF_X al_2e96e73a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[10]));
  AL_DFF_X al_48d21ce2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[11]));
  AL_DFF_X al_de16a3a5 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[12]));
  AL_DFF_X al_201c475f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[13]));
  AL_DFF_X al_13184e1c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_75776e99[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[0]));
  AL_DFF_X al_f302db52 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[1]));
  AL_DFF_X al_a80503f4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[2]));
  AL_DFF_X al_d897d548 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[3]));
  AL_DFF_X al_8e32cf6b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[4]));
  AL_DFF_X al_7b4e52a9 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[5]));
  AL_DFF_X al_215385fb (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[6]));
  AL_DFF_X al_b1daca73 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_bc5c8fc3[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(wave_sin[7]));
  AL_DFF_X al_ce6e5997 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[8]));
  AL_DFF_X al_7c322425 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[9]));
  AL_DFF_X al_1f65ec13 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[10]));
  AL_DFF_X al_5e904a35 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[0]));
  AL_DFF_X al_116f1db3 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[1]));
  AL_DFF_X al_6c993e82 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[2]));
  AL_DFF_X al_23963ea6 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[3]));
  AL_DFF_X al_6c25cf29 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[4]));
  AL_DFF_X al_e7cc423c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[5]));
  AL_DFF_X al_2c6ea385 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[6]));
  AL_DFF_X al_a356779f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8aaaf100[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6790cfef[7]));
  AL_DFF_X al_f27b108d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[8]));
  AL_DFF_X al_d1a67c2f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[9]));
  AL_DFF_X al_a7f95d18 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[10]));
  AL_DFF_X al_cbbb4490 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[0]));
  AL_DFF_X al_30153836 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[1]));
  AL_DFF_X al_37ead40d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[2]));
  AL_DFF_X al_7625712c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[3]));
  AL_DFF_X al_2531de5d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[4]));
  AL_DFF_X al_2ccbdc6d (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[5]));
  AL_DFF_X al_2c62c395 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[6]));
  AL_DFF_X al_ee1990ef (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_6790cfef[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8378b540[7]));
  AL_DFF_X al_db0079e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[8]));
  AL_DFF_X al_876f7db (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[9]));
  AL_DFF_X al_69a0ebce (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[10]));
  AL_DFF_X al_a6c89e95 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[11]));
  AL_DFF_X al_f3acd144 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[12]));
  AL_DFF_X al_e87e6f9a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_b33e7450[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[0]));
  AL_DFF_X al_43ae41e1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[1]));
  AL_DFF_X al_32098dc2 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[2]));
  AL_DFF_X al_1771790f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[3]));
  AL_DFF_X al_4e0fd4b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[4]));
  AL_DFF_X al_1d1fe749 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[5]));
  AL_DFF_X al_f8b279ec (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[6]));
  AL_DFF_X al_75a93bc1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_fcd55aa0[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_582c7f1a[7]));
  AL_DFF_X al_8117d99a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[8]));
  AL_DFF_X al_170fafe0 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[9]));
  AL_DFF_X al_d7229bc1 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[10]));
  AL_DFF_X al_d80ca115 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[11]));
  AL_DFF_X al_a73edca8 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[12]));
  AL_DFF_X al_2e8a2570 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[0]));
  AL_DFF_X al_4c05617e (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[1]));
  AL_DFF_X al_7cbb1b5f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[2]));
  AL_DFF_X al_1851373 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[3]));
  AL_DFF_X al_6ef4721c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[4]));
  AL_DFF_X al_ef14836c (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[5]));
  AL_DFF_X al_29111b42 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[6]));
  AL_DFF_X al_9e5c600b (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_defcae67[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cb3139[7]));
  AL_DFF_X al_8ff57d60 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[8]));
  AL_DFF_X al_47b511ab (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[9]));
  AL_DFF_X al_89005d1a (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[10]));
  AL_DFF_X al_f5b5ca38 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[11]));
  AL_DFF_X al_7907a48 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[12]));
  AL_DFF_X al_3176eb22 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_8378b540[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[0]));
  AL_DFF_X al_1ec04f80 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[1]));
  AL_DFF_X al_ec2280f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[2]));
  AL_DFF_X al_ecb5afd4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[3]));
  AL_DFF_X al_d15fb662 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[4]));
  AL_DFF_X al_e22992ea (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[5]));
  AL_DFF_X al_c3bb0c4f (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[6]));
  AL_DFF_X al_5b797485 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_d0d95c2b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c6da17f[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7b15ddba (
    .a(al_7cb3139[10]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[10]),
    .o(al_6b994b8c[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c82f5456 (
    .a(al_7cb3139[11]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[11]),
    .o(al_6b994b8c[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_9ce009e7 (
    .a(al_7cb3139[12]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[12]),
    .o(al_6b994b8c[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_367b458 (
    .a(al_8e2f713c),
    .b(al_cc82cb7d[13]),
    .o(al_6b994b8c[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c3b30651 (
    .a(al_7cb3139[1]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[1]),
    .o(al_6b994b8c[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_2b32cf8a (
    .a(al_7cb3139[2]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[2]),
    .o(al_6b994b8c[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_e2ac39fc (
    .a(al_7cb3139[3]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[3]),
    .o(al_6b994b8c[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_49ece604 (
    .a(al_7cb3139[4]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[4]),
    .o(al_6b994b8c[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_bef2872a (
    .a(al_7cb3139[5]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[5]),
    .o(al_6b994b8c[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_ebd5c0c4 (
    .a(al_7cb3139[6]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[6]),
    .o(al_6b994b8c[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_ab8f8a85 (
    .a(al_7cb3139[7]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[7]),
    .o(al_6b994b8c[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_465fe84 (
    .a(al_7cb3139[8]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[8]),
    .o(al_6b994b8c[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_55e58a6f (
    .a(al_7cb3139[9]),
    .b(al_8e2f713c),
    .c(al_cc82cb7d[9]),
    .o(al_6b994b8c[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_78e72845 (
    .a(al_411d7869[30]),
    .b(al_411d7869[31]),
    .o(al_5fbe7497));
  AL_DFF_X al_f27e26c4 (
    .ar(~rst_n),
    .as(1'b0),
    .clk(clk),
    .d(al_5fbe7497),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e2f713c));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d456667 (
    .a(al_75776e99[10]),
    .b(al_347def8c[31]),
    .c(al_747bea5[10]),
    .o(al_bc5c8fc3[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d9de8342 (
    .a(al_75776e99[11]),
    .b(al_347def8c[31]),
    .c(al_747bea5[11]),
    .o(al_bc5c8fc3[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c593df9f (
    .a(al_75776e99[12]),
    .b(al_347def8c[31]),
    .c(al_747bea5[12]),
    .o(al_bc5c8fc3[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fce59cb7 (
    .a(al_347def8c[31]),
    .b(al_747bea5[13]),
    .o(al_bc5c8fc3[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d6aba0b6 (
    .a(al_75776e99[1]),
    .b(al_347def8c[31]),
    .c(al_747bea5[1]),
    .o(al_bc5c8fc3[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_bba87de2 (
    .a(al_75776e99[2]),
    .b(al_347def8c[31]),
    .c(al_747bea5[2]),
    .o(al_bc5c8fc3[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a8d32043 (
    .a(al_75776e99[3]),
    .b(al_347def8c[31]),
    .c(al_747bea5[3]),
    .o(al_bc5c8fc3[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_c61147f4 (
    .a(al_75776e99[4]),
    .b(al_347def8c[31]),
    .c(al_747bea5[4]),
    .o(al_bc5c8fc3[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_b08d86be (
    .a(al_75776e99[5]),
    .b(al_347def8c[31]),
    .c(al_747bea5[5]),
    .o(al_bc5c8fc3[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_4326cc2d (
    .a(al_75776e99[6]),
    .b(al_347def8c[31]),
    .c(al_747bea5[6]),
    .o(al_bc5c8fc3[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_dfe3ec93 (
    .a(al_75776e99[7]),
    .b(al_347def8c[31]),
    .c(al_747bea5[7]),
    .o(al_bc5c8fc3[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_faff0718 (
    .a(al_75776e99[8]),
    .b(al_347def8c[31]),
    .c(al_747bea5[8]),
    .o(al_bc5c8fc3[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_249078a7 (
    .a(al_75776e99[9]),
    .b(al_347def8c[31]),
    .c(al_747bea5[9]),
    .o(al_bc5c8fc3[9]));

endmodule 

