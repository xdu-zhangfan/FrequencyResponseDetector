// Verilog netlist created by Tang Dynasty v5.6.71036
// Wed Jul 12 23:02:35 2023

`timescale 1ns / 1ps
module dds_divider_0
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [31:0] denominator;
  input [31:0] numerator;
  input rst;
  input start;
  output done;
  output [31:0] quotient;
  output [31:0] remainder;

  parameter PIPLE = 34;
  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 32;
  parameter W_NUM = 32;
  parameter W_REM = 32;
  // localparam INPUT_PIPLINE = 1'b1;
  // localparam ITERA_PIPLINE = 32'b11111111111111111111111111111111;
  // localparam OUTPUT_PIPLINE = 1'b1;
  // localparam SubSft[0].i = 0;
  // localparam SubSft[10].i = 10;
  // localparam SubSft[11].i = 11;
  // localparam SubSft[12].i = 12;
  // localparam SubSft[13].i = 13;
  // localparam SubSft[14].i = 14;
  // localparam SubSft[15].i = 15;
  // localparam SubSft[16].i = 16;
  // localparam SubSft[17].i = 17;
  // localparam SubSft[18].i = 18;
  // localparam SubSft[19].i = 19;
  // localparam SubSft[1].i = 1;
  // localparam SubSft[20].i = 20;
  // localparam SubSft[21].i = 21;
  // localparam SubSft[22].i = 22;
  // localparam SubSft[23].i = 23;
  // localparam SubSft[24].i = 24;
  // localparam SubSft[25].i = 25;
  // localparam SubSft[26].i = 26;
  // localparam SubSft[27].i = 27;
  // localparam SubSft[28].i = 28;
  // localparam SubSft[29].i = 29;
  // localparam SubSft[2].i = 2;
  // localparam SubSft[30].i = 30;
  // localparam SubSft[31].i = 31;
  // localparam SubSft[3].i = 3;
  // localparam SubSft[4].i = 4;
  // localparam SubSft[5].i = 5;
  // localparam SubSft[6].i = 6;
  // localparam SubSft[7].i = 7;
  // localparam SubSft[8].i = 8;
  // localparam SubSft[9].i = 9;
  wire [31:0] al_d3fd7d5a;
  wire [2:0] al_4b6a4daa;
  wire [52:0] al_6f9059d1;
  wire [31:0] al_f2b51288;
  wire [11:0] al_42afff14;
  wire [31:0] al_5d497694;
  wire [10:0] al_fac191b8;
  wire [2:0] al_adb04807;
  wire [51:0] al_177a13cd;
  wire [31:0] al_6c6869d7;
  wire [12:0] al_e45a58d8;
  wire [31:0] al_c2901510;
  wire [11:0] al_c9ed4b28;
  wire [2:0] al_2e1bd9dc;
  wire [50:0] al_a6f4a789;
  wire [31:0] al_13d2e70f;
  wire [13:0] al_39a3b856;
  wire [31:0] al_fb9cdc0e;
  wire [12:0] al_8fc8d46f;
  wire [2:0] al_c6d10c98;
  wire [49:0] al_515b933;
  wire [31:0] al_7cada4c1;
  wire [14:0] al_5ced65c5;
  wire [31:0] al_28d525d8;
  wire [13:0] al_a63aa325;
  wire [2:0] al_599810dd;
  wire [48:0] al_82ca84f8;
  wire [31:0] al_5fd65077;
  wire [15:0] al_51f816c9;
  wire [31:0] al_8d341179;
  wire [14:0] al_1898703d;
  wire [2:0] al_903e8807;
  wire [47:0] al_297c219f;
  wire [31:0] al_174c5039;
  wire [16:0] al_bcdd8ff0;
  wire [31:0] al_45052583;
  wire [15:0] al_ebfa785c;
  wire [2:0] al_5ed5f44b;
  wire [46:0] al_2e95330c;
  wire [31:0] al_1276f4f7;
  wire [17:0] al_d11b8;
  wire [31:0] al_b5df9b8a;
  wire [16:0] al_b4daf6f3;
  wire [2:0] al_54284e1f;
  wire [45:0] al_b4e2b23b;
  wire [31:0] al_3692f86e;
  wire [18:0] al_2bcf47f2;
  wire [31:0] al_28955387;
  wire [17:0] al_9c94ca47;
  wire [2:0] al_f83a6cd4;
  wire [44:0] al_e7d838f;
  wire [31:0] al_368cfa5b;
  wire [19:0] al_f57e3792;
  wire [31:0] al_e55e130b;
  wire [18:0] al_def6d145;
  wire [2:0] al_b0a2efb7;
  wire [43:0] al_30e951fe;
  wire [31:0] al_e240f99f;
  wire [20:0] al_755dcbd4;
  wire [31:0] al_abd7cd63;
  wire [19:0] al_bf1e6610;
  wire [2:0] al_3da4ff6f;
  wire [61:0] al_3bd314e4;
  wire [31:0] al_83a08f3f;
  wire [31:0] al_89f2771a;
  wire [1:0] al_33c3313d;
  wire [2:0] al_1c8da1e8;
  wire [42:0] al_e803eabe;
  wire [31:0] al_80a0f09e;
  wire [21:0] al_ceb4d3af;
  wire [31:0] al_cdad9264;
  wire [20:0] al_bd7f7f17;
  wire [2:0] al_acb3303d;
  wire [41:0] al_753f5f88;
  wire [31:0] al_98494645;
  wire [22:0] al_c706fd91;
  wire [31:0] al_f7ed724c;
  wire [21:0] al_be8c4478;
  wire [2:0] al_14a1a59a;
  wire [40:0] al_35594bd9;
  wire [31:0] al_bf34d64d;
  wire [23:0] al_abd8c6ec;
  wire [31:0] al_96533024;
  wire [22:0] al_f1d740ba;
  wire [2:0] al_21143207;
  wire [39:0] al_f2bb4ec4;
  wire [31:0] al_f0f43754;
  wire [24:0] al_801f6a4a;
  wire [31:0] al_e60d8647;
  wire [23:0] al_d3734717;
  wire [2:0] al_e0dc7e9e;
  wire [38:0] al_3029c49a;
  wire [31:0] al_86280a69;
  wire [25:0] al_591ecc80;
  wire [31:0] al_f78b30ce;
  wire [24:0] al_4a4fb8f1;
  wire [2:0] al_bade9fae;
  wire [37:0] al_5181785e;
  wire [31:0] al_9e3033a4;
  wire [26:0] al_b677b8b1;
  wire [31:0] al_63579c4c;
  wire [25:0] al_28f9bf01;
  wire [2:0] al_8f9ab06;
  wire [36:0] al_6a56028d;
  wire [31:0] al_7397600a;
  wire [27:0] al_64d71d5a;
  wire [31:0] al_2c297489;
  wire [26:0] al_c0ef3ebf;
  wire [2:0] al_fee4bd37;
  wire [35:0] al_b6768e55;
  wire [31:0] al_e4be4089;
  wire [28:0] al_c20bde66;
  wire [31:0] al_9857f6b5;
  wire [27:0] al_d71a2aba;
  wire [2:0] al_e0e2aae4;
  wire [34:0] al_222a5f4d;
  wire [31:0] al_4a463b38;
  wire [29:0] al_632b75dc;
  wire [31:0] al_e343d659;
  wire [28:0] al_c7a3cd65;
  wire [2:0] al_5db428bb;
  wire [33:0] al_d1a07609;
  wire [31:0] al_32ba5b24;
  wire [30:0] al_10f8c714;
  wire [31:0] al_14165a56;
  wire [29:0] al_bad3f013;
  wire [2:0] al_67f5b0b3;
  wire [60:0] al_6a637a32;
  wire [31:0] al_3d0cfeb4;
  wire [31:0] al_a9b28455;
  wire [2:0] al_b54c1014;
  wire [2:0] al_8d805738;
  wire [32:0] al_627988c3;
  wire [31:0] al_690b21a4;
  wire [31:0] al_7c1783ce;
  wire [31:0] al_3ccb3a4f;
  wire [30:0] al_9d67405f;
  wire [2:0] al_74993dd2;
  wire [31:0] al_a5e9c08d;
  wire [31:0] al_57dc9b0c;
  wire [31:0] al_eb7d14b9;
  wire [32:0] al_df3b43b5;
  wire [31:0] al_b40233aa;
  wire [2:0] al_44882eca;
  wire [59:0] al_b052c226;
  wire [31:0] al_592f1b09;
  wire [4:0] al_828cf6c5;
  wire [31:0] al_8c015879;
  wire [3:0] al_b18b7cbb;
  wire [2:0] al_f336c405;
  wire [58:0] al_28202fa7;
  wire [31:0] al_1d4399b1;
  wire [31:0] al_7a8c14f1;
  wire [4:0] al_917df14b;
  wire [2:0] al_f23786d8;
  wire [57:0] al_68bb3ebd;
  wire [31:0] al_1b3e91c5;
  wire [6:0] al_d01f30c3;
  wire [31:0] al_7d7cdb8e;
  wire [5:0] al_4682e2e2;
  wire [2:0] al_6e4d5f5f;
  wire [56:0] al_f2a9de02;
  wire [31:0] al_15503509;
  wire [7:0] al_f3dd9213;
  wire [31:0] al_78306f09;
  wire [6:0] al_22a22ff3;
  wire [2:0] al_d255f877;
  wire [55:0] al_5206392b;
  wire [31:0] al_59bef53b;
  wire [8:0] al_727f921;
  wire [31:0] al_601b9c02;
  wire [7:0] al_9c3e2402;
  wire [2:0] al_30922aac;
  wire [54:0] al_d6cb04b6;
  wire [31:0] al_f7a9a92b;
  wire [9:0] al_96e7074d;
  wire [31:0] al_3b7f0416;
  wire [8:0] al_4dd3fb65;
  wire [2:0] al_36d845bb;
  wire [53:0] al_c1960abd;
  wire [31:0] al_5283b07c;
  wire [10:0] al_c855b680;
  wire [31:0] al_bcaebe78;
  wire [9:0] al_3cd0a9ea;
  wire [2:0] al_ae5d831a;
  wire [62:0] al_9d1d5c0;
  wire [31:0] al_a5806bc7;
  wire [31:0] al_3519ff8d;
  wire [31:0] al_18157fe8;
  wire al_51794c84;
  wire al_8d24c5a7;
  wire al_bff2070;
  wire al_d6a2c880;
  wire al_25015351;
  wire al_a11c1e55;
  wire al_7cfee86d;
  wire al_b80fa848;
  wire al_9bab634c;
  wire al_c65e897c;
  wire al_428c242;
  wire al_5aafa5e1;
  wire al_d2131a9e;
  wire al_67364858;
  wire al_d83723e4;
  wire al_493db12b;
  wire al_d6eab53e;
  wire al_dfe53854;
  wire al_b97fef0c;
  wire al_ee38d1b0;
  wire al_bbc0fba0;
  wire al_e8cc505e;
  wire al_9f82cc8e;
  wire al_784f99f2;
  wire al_818d701;
  wire al_b3f0117a;
  wire al_e3a4cb77;
  wire al_6c8e3937;
  wire al_dbc3e2b0;
  wire al_a04b98a0;
  wire al_e0aedfd3;
  wire al_150d105b;
  wire al_6f78cae7;
  wire al_2e62154a;
  wire al_e5b9a180;
  wire al_a4e131c6;
  wire al_7087d50d;
  wire al_6b08641e;
  wire al_b95fb7ea;
  wire al_ac18f4f8;
  wire al_8cbaef5d;
  wire al_8c892fd7;
  wire al_eb1649fe;
  wire al_7b45fe04;
  wire al_8035eade;
  wire al_42e0e24e;
  wire al_71245cc2;
  wire al_32780627;
  wire al_65eed942;
  wire al_74dcac58;
  wire al_5da4a00d;
  wire al_beb32d78;
  wire al_32d68c1d;
  wire al_41f22393;
  wire al_28817105;
  wire al_93c58a47;
  wire al_8b10921e;
  wire al_806ca727;
  wire al_f4ebe63d;
  wire al_b1ae99ca;
  wire al_c7b36065;
  wire al_466d66e9;
  wire al_cb6f9733;
  wire al_884856d;
  wire al_d72d321f;
  wire al_5742b37b;
  wire al_e4c6cc49;
  wire al_6f18daeb;
  wire al_3fd86060;
  wire al_7fd69b02;
  wire al_3b5f5572;
  wire al_926f19c9;
  wire al_71819c0f;
  wire al_16cd5903;
  wire al_f4b0959f;
  wire al_b87d9ba8;
  wire al_415da9aa;
  wire al_8465c727;
  wire al_f7c19df7;
  wire al_3ed120c9;
  wire al_3f4489bf;
  wire al_ae5b1fc6;
  wire al_858ee963;
  wire al_c2097ceb;
  wire al_1f755058;
  wire al_1c729801;
  wire al_cc2d4a37;
  wire al_171301db;
  wire al_b8a0b712;
  wire al_5c73d821;
  wire al_6d30b4d3;
  wire al_c8e591e5;
  wire al_ba0cc25;
  wire al_3df74a2f;
  wire al_2265cd1e;
  wire al_eeaf7eee;
  wire al_99a412d5;
  wire al_6fc7ef08;
  wire al_60f2f1ac;
  wire al_fbd5879f;
  wire al_1800fb32;
  wire al_6bb8dfe8;
  wire al_a8cd8f3c;
  wire al_d4a26700;
  wire al_632a2e97;
  wire al_6222dcd7;
  wire al_78a5b5c9;
  wire al_9eeae501;
  wire al_c05929c6;
  wire al_b2191d5e;
  wire al_f7339674;
  wire al_6ded130e;
  wire al_467f742e;
  wire al_1cf1391b;
  wire al_d649f6ed;
  wire al_d568756b;
  wire al_3f5f9369;
  wire al_cad8537e;
  wire al_def1a789;
  wire al_e869e5fb;
  wire al_38880c22;
  wire al_74d32fe0;
  wire al_f930adec;
  wire al_3cd6c50e;
  wire al_d4f61208;
  wire al_cc07f579;
  wire al_9d3c2203;
  wire al_c3c604b3;
  wire al_949714ad;
  wire al_691c6b01;
  wire al_aa40ea6e;
  wire al_dad76b0c;
  wire al_a0c202f4;
  wire al_3ec72efd;
  wire al_64c5377c;
  wire al_499f819a;
  wire al_d3b6fe74;
  wire al_efcf8b1a;
  wire al_e9939d22;
  wire al_b2bc9399;
  wire al_96577a6c;
  wire al_a511a420;
  wire al_523c4f95;
  wire al_be2eadc2;
  wire al_1bf3430d;
  wire al_ee8cd800;
  wire al_289b6994;
  wire al_278e8e9c;
  wire al_62d4794d;
  wire al_9d67c14b;
  wire al_5d2d77b4;
  wire al_37d85dd8;
  wire al_22c0f879;
  wire al_a6323dfd;
  wire al_d459fd2a;
  wire al_a0f8478c;
  wire al_67dd1cc2;
  wire al_9380c67b;
  wire al_6b7d50a7;
  wire al_4cc7f121;
  wire al_648c2518;
  wire al_1ba5074a;
  wire al_959737fa;
  wire al_456e9f5b;
  wire al_983289c4;
  wire al_170bfe43;
  wire al_96c24183;
  wire al_a7a2d586;
  wire al_1ba7203c;
  wire al_fdbea65d;
  wire al_92ca20ed;
  wire al_2758bb5;
  wire al_337113ba;
  wire al_579fe9c9;
  wire al_b98fe565;
  wire al_60ed0a3f;
  wire al_27d9400d;
  wire al_94badae1;
  wire al_462fcfec;
  wire al_11444b05;
  wire al_6a490a84;
  wire al_7c4effa7;
  wire al_2a54b225;
  wire al_bf2e29ab;
  wire al_1741bada;
  wire al_506041c3;
  wire al_ff00a5b;
  wire al_cadab979;
  wire al_1ca453a8;
  wire al_a7dd3d61;
  wire al_f0c84e95;
  wire al_11666a8e;
  wire al_2f88a0b8;
  wire al_6a534ff7;
  wire al_22cba5b6;
  wire al_dc8a8f4;
  wire al_3ad2f5fe;
  wire al_877d1bc;
  wire al_80347035;
  wire al_54975822;
  wire al_e5f75e51;
  wire al_84743aea;
  wire al_4c6c1136;
  wire al_aff6af71;
  wire al_786cd6fa;
  wire al_ea94f7fb;
  wire al_83614d40;
  wire al_4182734;
  wire al_c006efbd;
  wire al_49456793;
  wire al_e7a93f78;
  wire al_dd519345;
  wire al_842cba6d;
  wire al_bf0c2f5d;
  wire al_5059c5b1;
  wire al_cf4d3fd;
  wire al_1df89094;
  wire al_fdd90390;
  wire al_6e7e6fcf;
  wire al_2daedad1;
  wire al_3b13cff4;
  wire al_cc19a77c;
  wire al_e8916352;
  wire al_3317fa82;
  wire al_2ca9607b;
  wire al_90792e1b;
  wire al_2af03fa4;
  wire al_9b8ff49a;
  wire al_b2d82920;
  wire al_13bec3a1;
  wire al_62013390;
  wire al_885349b2;
  wire al_905b8225;
  wire al_ebf67b92;
  wire al_e856fef8;
  wire al_3b01c73c;
  wire al_5f9be50;
  wire al_c495520b;
  wire al_31fa6069;
  wire al_add99006;
  wire al_3c7582f0;
  wire al_ad366bd4;
  wire al_435dca9c;
  wire al_5689e405;
  wire al_af9115e4;
  wire al_60435cbc;
  wire al_e0c9a948;
  wire al_402ba912;
  wire al_8caee7aa;
  wire al_b7e03ff;
  wire al_74039666;
  wire al_9da6bf97;
  wire al_23c46bef;
  wire al_8c81e3ca;
  wire al_f64316;
  wire al_be55634f;
  wire al_631a2483;
  wire al_f8dbc1a1;
  wire al_ba13973b;
  wire al_e67fe640;
  wire al_7f8fdeae;
  wire al_9d447f48;
  wire al_56164bd3;
  wire al_f9511aee;
  wire al_6a25f3ea;
  wire al_abf34df7;
  wire al_a6796ab;
  wire al_59ba0f55;
  wire al_92ed39a9;
  wire al_c6dcc95e;
  wire al_1f87453b;
  wire al_4c52cca8;
  wire al_bf05760;
  wire al_ceb7552e;
  wire al_56dc547b;
  wire al_cd3ff18;
  wire al_cee7ade2;
  wire al_afdea3b6;
  wire al_ed22eb5b;
  wire al_7894a2ed;
  wire al_c319c1b9;
  wire al_3111d364;
  wire al_4e50336d;
  wire al_99511a1d;
  wire al_c83520d8;
  wire al_d6fc0fa3;
  wire al_5b46bf26;
  wire al_5094d9fc;
  wire al_94cd1325;
  wire al_b9861408;
  wire al_976c5f9d;
  wire al_e586ffc9;
  wire al_b45c14e1;
  wire al_1b1dea64;
  wire al_4188fe4e;
  wire al_de74a82;
  wire al_632e424b;
  wire al_7fd8d148;
  wire al_6d674526;
  wire al_fdad78c8;
  wire al_6620847d;
  wire al_f4867e16;
  wire al_1bdf229b;
  wire al_3e7ed8c8;
  wire al_354fda56;
  wire al_2f8d1c1e;
  wire al_57929d06;
  wire al_325baf0c;
  wire al_9079498a;
  wire al_d2dbac27;
  wire al_7715910d;
  wire al_f486a09d;
  wire al_bee033d9;
  wire al_a60df36b;
  wire al_aa119f92;
  wire al_ced042bc;
  wire al_9de12621;
  wire al_c6d35f30;
  wire al_41de2ced;
  wire al_a4baa375;
  wire al_7d7301fd;
  wire al_f804f442;
  wire al_fa20e924;
  wire al_75df31c;
  wire al_fb6c6a88;
  wire al_6a47eaf1;
  wire al_ef2cb93b;
  wire al_7c6e81bc;
  wire al_820ba18b;
  wire al_90eca21f;
  wire al_14135fe;
  wire al_278fc7b9;
  wire al_78f968d6;
  wire al_6cb6cc70;
  wire al_5bfcf8ca;
  wire al_7777e58e;
  wire al_ce2d0e53;
  wire al_665b7858;
  wire al_3d0d887e;
  wire al_f44c949b;
  wire al_394ce23b;
  wire al_354fae1f;
  wire al_89af750e;
  wire al_8cf6cbd4;
  wire al_32030ed2;
  wire al_5875f740;
  wire al_7cb5ff51;
  wire al_ee0cbe48;
  wire al_b4749ad8;
  wire al_dc8ef999;
  wire al_500654bb;
  wire al_62272aaf;
  wire al_2f455704;
  wire al_b7b82cb6;
  wire al_7375cfb0;
  wire al_c78e76e7;
  wire al_ef33e959;
  wire al_6387fe;
  wire al_25d9aae7;
  wire al_9233bdf0;
  wire al_cee8b982;
  wire al_c5ec6219;
  wire al_ae24ecf8;
  wire al_72ba4be2;
  wire al_3a745b61;
  wire al_2878e2ee;
  wire al_1abbaba6;
  wire al_ec19d56e;
  wire al_6409430b;
  wire al_33374be5;
  wire al_97f76d83;
  wire al_111f57ad;
  wire al_dd5d3b13;
  wire al_daa9922c;
  wire al_d0a99602;
  wire al_5a02bf80;
  wire al_67d1c21c;
  wire al_e79544d1;
  wire al_8f3b225e;
  wire al_b10d3e54;
  wire al_fa88be3f;
  wire al_17625a21;
  wire al_19e00ab1;
  wire al_c7f6f4df;
  wire al_ea4ffb3c;
  wire al_e688eccb;
  wire al_ec10f532;
  wire al_a1afdc44;
  wire al_d4e70d9d;
  wire al_16d28d90;
  wire al_48808c89;
  wire al_6216f648;
  wire al_71a4da9;
  wire al_f45fae5e;
  wire al_d7aedbc5;
  wire al_754bf737;
  wire al_7fd7f68e;
  wire al_b3ed3b7d;
  wire al_c41f5a7c;
  wire al_f31b3480;
  wire al_864bc6dc;
  wire al_f693e61d;
  wire al_47955db6;
  wire al_cc078df4;
  wire al_58dab36d;
  wire al_3e035452;
  wire al_106a827;
  wire al_f709c5ab;
  wire al_56abe384;
  wire al_7418c94f;
  wire al_efa49dac;
  wire al_e130ad23;
  wire al_2f299606;
  wire al_925eb901;
  wire al_daeef93a;
  wire al_2ff932f4;
  wire al_2e6e4c5b;
  wire al_2a6886e2;
  wire al_1f220fb;
  wire al_7154b9a7;
  wire al_1bf81a9b;
  wire al_1b451831;
  wire al_72e17b7c;
  wire al_a1fc4ea8;
  wire al_dde82c43;
  wire al_b1d329d9;
  wire al_c8aee28f;
  wire al_b33e7544;
  wire al_accca793;
  wire al_4dd25e15;
  wire al_c76b4c37;
  wire al_b7a54e24;
  wire al_85587067;
  wire al_1ff06f87;
  wire al_143fe859;
  wire al_cd6d2794;
  wire al_e59fc5bd;
  wire al_bd4c5933;
  wire al_6c260918;
  wire al_6b532b61;
  wire al_9cdbacea;
  wire al_232548;
  wire al_e1d75325;
  wire al_87178f5;
  wire al_70012e88;
  wire al_452820cd;
  wire al_392bc465;
  wire al_adc3cec6;
  wire al_852fa027;
  wire al_3c9f5595;
  wire al_829de986;
  wire al_e3bf1d53;
  wire al_e6964d98;
  wire al_188e472a;
  wire al_d8b8a6e2;
  wire al_8044404c;
  wire al_ca8e61e8;
  wire al_3144b627;
  wire al_cb5d4eb2;
  wire al_e2af005f;
  wire al_dd8f16d1;
  wire al_f2a22ed1;
  wire al_d1a88ad2;
  wire al_3c316ef;
  wire al_a2fff3ec;
  wire al_f6ffe199;
  wire al_aa4c6187;
  wire al_3d105014;
  wire al_f0daa0db;
  wire al_47c0210d;
  wire al_85b1bb55;
  wire al_ebd1e7fe;
  wire al_bc14fb86;
  wire al_dd5db619;
  wire al_3e3b2341;
  wire al_9b3654ad;
  wire al_100303d6;
  wire al_50e17485;
  wire al_3b8d6cb9;
  wire al_83167981;
  wire al_3fb5c0bf;
  wire al_f7a0a5e;
  wire al_28c3840c;
  wire al_a5df252b;
  wire al_855effe8;
  wire al_966d3a1d;
  wire al_f4c9a2d4;
  wire al_42dadf79;
  wire al_97bfe275;
  wire al_8ef4e9d1;
  wire al_1a4fdc2c;
  wire al_99c43840;
  wire al_98c65d85;
  wire al_5b6cf04f;
  wire al_ae08306c;
  wire al_7f4546cf;
  wire al_f23b4ac3;
  wire al_ac9e4212;
  wire al_78275fb6;
  wire al_9a080fbf;
  wire al_8a23505f;
  wire al_5f9068e6;
  wire al_a46f14d2;
  wire al_342b0ff9;
  wire al_e782992a;
  wire al_5d589bca;
  wire al_33f64520;
  wire al_e9c34253;
  wire al_d36ef0a6;
  wire al_dd36b780;
  wire al_232ecfaf;
  wire al_f2fd9563;
  wire al_4c3e9ef3;
  wire al_6c944eaa;
  wire al_8f677fc9;
  wire al_5fcd8d3b;
  wire al_5fd9abe8;
  wire al_6c21e4f;
  wire al_1a0f9e95;
  wire al_56a083ea;
  wire al_7028725;
  wire al_aa188274;
  wire al_78d777d2;
  wire al_6769a627;
  wire al_249d4728;
  wire al_853654c1;
  wire al_5173861b;
  wire al_7a77d617;
  wire al_4f5a23d4;
  wire al_3eebd40f;
  wire al_8e4361ca;
  wire al_912de09d;
  wire al_85cca751;
  wire al_ad8d6e84;
  wire al_5992e66f;
  wire al_53645fd3;
  wire al_5c00f664;
  wire al_a5fb5d66;
  wire al_bfb57bee;
  wire al_2f85c10c;
  wire al_ce21f8f3;
  wire al_83736e7b;
  wire al_c3f591aa;
  wire al_fbb0bdd6;
  wire al_eb11562b;
  wire al_15d2d0ed;
  wire al_a792d40a;
  wire al_92024dcf;
  wire al_60518bd5;
  wire al_a0662365;
  wire al_d44591b2;
  wire al_1280dac2;
  wire al_655899d3;
  wire al_3a98aee3;
  wire al_6269677;
  wire al_f6aa030f;
  wire al_1e3baa15;
  wire al_90c4774;
  wire al_2d7cd5be;
  wire al_41002c4f;
  wire al_b06c909;
  wire al_bb31a1fd;
  wire al_52f7b6db;
  wire al_a8fa8fea;
  wire al_b2ffd084;
  wire al_b701d480;
  wire al_97262af6;
  wire al_2a480b9e;
  wire al_d720b206;
  wire al_b05ac301;
  wire al_67046fd1;
  wire al_108156ff;
  wire al_162e0df5;
  wire al_61845f15;
  wire al_17de8af8;
  wire al_e9f8df12;
  wire al_e7a7f7d2;
  wire al_37282f35;
  wire al_e1b1cb21;
  wire al_eb87db38;
  wire al_8db59e87;
  wire al_8fa4d3c;
  wire al_eddac2b0;
  wire al_a23f6f13;
  wire al_52cd72b8;
  wire al_a35c5ad0;
  wire al_bf78ad38;
  wire al_f71c0797;
  wire al_2d1a2942;
  wire al_c045eda5;
  wire al_892befbc;
  wire al_19974a3;
  wire al_634f8236;
  wire al_f607f1c2;
  wire al_42f85898;
  wire al_7269924;
  wire al_54056c79;
  wire al_3b37ef98;
  wire al_d63c55c7;
  wire al_dc0ce6da;
  wire al_8691ef65;
  wire al_ecc3713;
  wire al_de5112e6;
  wire al_6c82a93e;
  wire al_4a1ebbca;
  wire al_9535661e;
  wire al_90a06cdf;
  wire al_4f7fb1ad;
  wire al_f96974bd;
  wire al_6f00a1da;
  wire al_2f03a26;
  wire al_82784f18;
  wire al_2281381d;
  wire al_1e591849;
  wire al_e40698dd;
  wire al_552d5319;
  wire al_cadea4c8;
  wire al_203d257f;
  wire al_ca8f2e4c;
  wire al_ed33bb97;
  wire al_2be1d9b7;
  wire al_57ac52e7;
  wire al_5f980ce9;
  wire al_a2de35e1;
  wire al_4ba9ed11;
  wire al_cacb9d80;
  wire al_1bad0a7d;
  wire al_58234d6b;
  wire al_c5f2b310;
  wire al_477c87;
  wire al_b103a97e;
  wire al_d405f4db;
  wire al_59bc69f9;
  wire al_cb5c1242;
  wire al_b8df04a0;
  wire al_93714d98;
  wire al_f3cdefe2;
  wire al_25f6edd0;
  wire al_4b9b0b4;
  wire al_4ecce1a8;
  wire al_a74a382d;
  wire al_fa0c3c8b;
  wire al_67ed9c11;
  wire al_f563230a;
  wire al_c539d3e8;
  wire al_79960e7c;
  wire al_a9fdceb9;
  wire al_c9a744c1;
  wire al_631391e1;
  wire al_126d5412;
  wire al_7c9dcdbf;
  wire al_4de4f552;
  wire al_753472e;
  wire al_15e33bf2;
  wire al_64c930a8;
  wire al_6ff407e;
  wire al_ff0e3144;
  wire al_f8599920;
  wire al_b9af15ec;
  wire al_47c20a17;
  wire al_f5506553;
  wire al_a989c55e;
  wire al_6dfedbe6;
  wire al_cce5b1fa;
  wire al_682ed5c4;
  wire al_75a022;
  wire al_81b3dbd9;
  wire al_1fc14639;
  wire al_d1df1e3c;
  wire al_c46bddb5;
  wire al_24bfc94c;
  wire al_92dd4899;
  wire al_79a8092a;
  wire al_7e098907;
  wire al_ad4f86b8;
  wire al_a5ca0ead;
  wire al_ef88efba;
  wire al_15966972;
  wire al_75ca1e75;
  wire al_f0189703;
  wire al_9fc9935f;
  wire al_b37de4b4;
  wire al_7eb6704d;
  wire al_4d58224c;
  wire al_d150e9d;
  wire al_be714bda;
  wire al_62b2844e;
  wire al_23344b64;
  wire al_aa529150;
  wire al_d6b6abb7;
  wire al_7cd30609;
  wire al_9765a29c;
  wire al_9d15fc0c;
  wire al_8fcf5341;
  wire al_5e79a92a;
  wire al_8fff10ae;
  wire al_bf66278b;
  wire al_ec79a3f9;
  wire al_b02d6cd0;
  wire al_c5e93959;
  wire al_dfb70c9;
  wire al_f058aa98;

  AL_MAP_LUT6 #(
    .EQN("(D*C*B*A*~(~F*E))"),
    .INIT(64'h8000800000008000))
    al_9dff2df0 (
    .a(al_d6a2c880),
    .b(al_a11c1e55),
    .c(al_7cfee86d),
    .d(al_b80fa848),
    .e(al_9d1d5c0[31]),
    .f(al_a5806bc7[31]),
    .o(al_9bab634c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_26cf0d17 (
    .a(al_9d1d5c0[42]),
    .b(al_9d1d5c0[43]),
    .c(al_9d1d5c0[44]),
    .d(al_9d1d5c0[45]),
    .e(al_9d1d5c0[46]),
    .f(al_9d1d5c0[47]),
    .o(al_8d24c5a7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1a5436e8 (
    .a(al_9d1d5c0[36]),
    .b(al_9d1d5c0[37]),
    .c(al_9d1d5c0[38]),
    .d(al_9d1d5c0[39]),
    .e(al_9d1d5c0[40]),
    .f(al_9d1d5c0[41]),
    .o(al_7cfee86d));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_9b4706c1 (
    .a(al_9d1d5c0[32]),
    .b(al_9d1d5c0[33]),
    .c(al_9d1d5c0[34]),
    .d(al_9d1d5c0[35]),
    .e(al_9d1d5c0[62]),
    .o(al_b80fa848));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E*D*C*B*A))"),
    .INIT(64'h7fffffff00000000))
    al_484a2a84 (
    .a(al_d6a2c880),
    .b(al_a11c1e55),
    .c(al_7cfee86d),
    .d(al_b80fa848),
    .e(al_9d1d5c0[31]),
    .f(al_a5806bc7[31]),
    .o(al_d3fd7d5a[31]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_a8379a88 (
    .a(al_9d1d5c0[58]),
    .b(al_9d1d5c0[59]),
    .c(al_9d1d5c0[60]),
    .d(al_9d1d5c0[61]),
    .o(al_bff2070));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_5b25dce5 (
    .a(al_8d24c5a7),
    .b(al_bff2070),
    .c(al_9d1d5c0[56]),
    .d(al_9d1d5c0[57]),
    .o(al_d6a2c880));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_f4a16149 (
    .a(al_9d1d5c0[52]),
    .b(al_9d1d5c0[53]),
    .c(al_9d1d5c0[54]),
    .d(al_9d1d5c0[55]),
    .o(al_25015351));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_e456193d (
    .a(al_25015351),
    .b(al_9d1d5c0[48]),
    .c(al_9d1d5c0[49]),
    .d(al_9d1d5c0[50]),
    .e(al_9d1d5c0[51]),
    .o(al_a11c1e55));
  AL_DFF_X al_8dce07d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_51794c84),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3da4ff6f[0]));
  AL_DFF_X al_f17869c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[30]));
  AL_DFF_X al_6fdc1f90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[31]));
  AL_DFF_X al_44d9ad93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[32]));
  AL_DFF_X al_679776b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[33]));
  AL_DFF_X al_387e2ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[34]));
  AL_DFF_X al_80a1b5c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[35]));
  AL_DFF_X al_82721c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[36]));
  AL_DFF_X al_a3d5903 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[37]));
  AL_DFF_X al_e592a0e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[38]));
  AL_DFF_X al_acbeffc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[39]));
  AL_DFF_X al_4489e3a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[40]));
  AL_DFF_X al_d24980be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[41]));
  AL_DFF_X al_19345fce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[42]));
  AL_DFF_X al_a83a1d68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[43]));
  AL_DFF_X al_4e415d95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[44]));
  AL_DFF_X al_e9d17faf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[45]));
  AL_DFF_X al_f9de33b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[46]));
  AL_DFF_X al_9eaed2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[47]));
  AL_DFF_X al_b9ea836d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[48]));
  AL_DFF_X al_7b1dc668 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[49]));
  AL_DFF_X al_94e1ec6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[50]));
  AL_DFF_X al_62750b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[51]));
  AL_DFF_X al_d5e4ced0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[52]));
  AL_DFF_X al_f52612fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[53]));
  AL_DFF_X al_3bc1f989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[54]));
  AL_DFF_X al_6c2255e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[55]));
  AL_DFF_X al_86cc6f60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[56]));
  AL_DFF_X al_6eeb6b45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[57]));
  AL_DFF_X al_7e9e25ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[58]));
  AL_DFF_X al_87e3e56e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[59]));
  AL_DFF_X al_1039c870 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[60]));
  AL_DFF_X al_31609b5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[61]));
  AL_DFF_X al_3e667d37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[8]));
  AL_DFF_X al_76077a7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[9]));
  AL_DFF_X al_ca2bda3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[10]));
  AL_DFF_X al_aedcb3d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[11]));
  AL_DFF_X al_ddbd2522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[12]));
  AL_DFF_X al_eb7451b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[13]));
  AL_DFF_X al_1a5403e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[14]));
  AL_DFF_X al_aba09c80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[15]));
  AL_DFF_X al_3555f910 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[16]));
  AL_DFF_X al_6cf7f1dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[17]));
  AL_DFF_X al_303c087 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[0]));
  AL_DFF_X al_be5dd8e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[18]));
  AL_DFF_X al_337785ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[19]));
  AL_DFF_X al_40b69221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[20]));
  AL_DFF_X al_a0f33db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[21]));
  AL_DFF_X al_556bbfeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[22]));
  AL_DFF_X al_98431931 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[23]));
  AL_DFF_X al_4bd4ce05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[24]));
  AL_DFF_X al_b17b5a51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[25]));
  AL_DFF_X al_149ddc26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[26]));
  AL_DFF_X al_21d87ca5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[27]));
  AL_DFF_X al_111950cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[1]));
  AL_DFF_X al_e9561921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[28]));
  AL_DFF_X al_a32c087c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[29]));
  AL_DFF_X al_7ebb2209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[30]));
  AL_DFF_X al_f66eda48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3fd7d5a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[31]));
  AL_DFF_X al_2f2000a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[2]));
  AL_DFF_X al_55e6c491 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[3]));
  AL_DFF_X al_d8753092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[4]));
  AL_DFF_X al_d994f8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[5]));
  AL_DFF_X al_cda80bef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[6]));
  AL_DFF_X al_da8e3c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[7]));
  AL_DFF_X al_b01a1a07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bab634c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33c3313d[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7275908b (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .o(al_e3a4cb77));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_289aaade (
    .a(1'b0),
    .o({al_c65e897c,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d6a2f7f9 (
    .a(al_f2b51288[21]),
    .b(al_6f9059d1[21]),
    .c(al_c65e897c),
    .o({al_428c242,al_42afff14[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7ab18fd (
    .a(al_f2b51288[22]),
    .b(al_6f9059d1[22]),
    .c(al_428c242),
    .o({al_5aafa5e1,al_42afff14[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed749a90 (
    .a(al_f2b51288[23]),
    .b(al_6f9059d1[23]),
    .c(al_5aafa5e1),
    .o({al_d2131a9e,al_42afff14[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_46115c4c (
    .a(al_f2b51288[24]),
    .b(al_6f9059d1[24]),
    .c(al_d2131a9e),
    .o({al_67364858,al_42afff14[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_776d0cd0 (
    .a(al_f2b51288[25]),
    .b(al_6f9059d1[25]),
    .c(al_67364858),
    .o({al_d83723e4,al_42afff14[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6eb8f4c (
    .a(al_f2b51288[26]),
    .b(al_6f9059d1[26]),
    .c(al_d83723e4),
    .o({al_493db12b,al_42afff14[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f2a100b (
    .a(al_f2b51288[27]),
    .b(al_6f9059d1[27]),
    .c(al_493db12b),
    .o({al_d6eab53e,al_42afff14[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33f1713e (
    .a(al_f2b51288[28]),
    .b(al_6f9059d1[28]),
    .c(al_d6eab53e),
    .o({al_dfe53854,al_42afff14[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a809cdcc (
    .a(al_f2b51288[29]),
    .b(al_6f9059d1[29]),
    .c(al_dfe53854),
    .o({al_b97fef0c,al_42afff14[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b31cc59e (
    .a(al_f2b51288[30]),
    .b(al_6f9059d1[30]),
    .c(al_b97fef0c),
    .o({al_ee38d1b0,al_42afff14[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ff01b79 (
    .a(al_f2b51288[31]),
    .b(al_6f9059d1[31]),
    .c(al_ee38d1b0),
    .o({al_bbc0fba0,al_42afff14[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a556e0b (
    .c(al_bbc0fba0),
    .o({open_n5,al_42afff14[11]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1017b365 (
    .a(al_6f9059d1[35]),
    .b(al_6f9059d1[36]),
    .c(al_6f9059d1[37]),
    .d(al_6f9059d1[38]),
    .e(al_6f9059d1[39]),
    .f(al_6f9059d1[40]),
    .o(al_e8cc505e));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_a98c8e1 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[0]),
    .e(al_f2b51288[21]),
    .o(al_5d497694[21]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_96b45486 (
    .a(al_6f9059d1[43]),
    .b(al_6f9059d1[44]),
    .c(al_6f9059d1[45]),
    .d(al_6f9059d1[46]),
    .o(al_9f82cc8e));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_c186dabe (
    .a(al_e8cc505e),
    .b(al_9f82cc8e),
    .c(al_6f9059d1[41]),
    .d(al_6f9059d1[42]),
    .o(al_784f99f2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_dd8ba473 (
    .a(al_6f9059d1[47]),
    .b(al_6f9059d1[48]),
    .c(al_6f9059d1[49]),
    .d(al_6f9059d1[50]),
    .e(al_6f9059d1[51]),
    .f(al_6f9059d1[52]),
    .o(al_818d701));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_92dfaa16 (
    .a(al_42afff14[11]),
    .b(al_6f9059d1[32]),
    .c(al_6f9059d1[33]),
    .d(al_6f9059d1[34]),
    .o(al_b3f0117a));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_180e0843 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[1]),
    .e(al_f2b51288[22]),
    .o(al_5d497694[22]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_4f03d1d (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[2]),
    .e(al_f2b51288[23]),
    .o(al_5d497694[23]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_9eee7f5b (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[3]),
    .e(al_f2b51288[24]),
    .o(al_5d497694[24]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_72963483 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[4]),
    .e(al_f2b51288[25]),
    .o(al_5d497694[25]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_798d52ce (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[5]),
    .e(al_f2b51288[26]),
    .o(al_5d497694[26]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_965ee5e8 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[6]),
    .e(al_f2b51288[27]),
    .o(al_5d497694[27]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_7f4b6f41 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[7]),
    .e(al_f2b51288[28]),
    .o(al_5d497694[28]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_a55b3215 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[8]),
    .e(al_f2b51288[29]),
    .o(al_5d497694[29]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_edf6097d (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[9]),
    .e(al_f2b51288[30]),
    .o(al_5d497694[30]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((C*B*A))+E*D*~((C*B*A))+~(E)*D*(C*B*A)+E*D*(C*B*A))"),
    .INIT(32'hff7f8000))
    al_6a52b4b9 (
    .a(al_784f99f2),
    .b(al_818d701),
    .c(al_b3f0117a),
    .d(al_42afff14[10]),
    .e(al_f2b51288[31]),
    .o(al_5d497694[31]));
  AL_DFF_X al_b4281495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4b6a4daa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adb04807[0]));
  AL_DFF_X al_cbebd2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[20]));
  AL_DFF_X al_a8473def (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[21]));
  AL_DFF_X al_c468c4fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[22]));
  AL_DFF_X al_e54f4c66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[23]));
  AL_DFF_X al_c371e0fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[24]));
  AL_DFF_X al_b0ef233c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[25]));
  AL_DFF_X al_582ed9cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[26]));
  AL_DFF_X al_df82421e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[27]));
  AL_DFF_X al_8cd4c4d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[28]));
  AL_DFF_X al_4e479f51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[29]));
  AL_DFF_X al_5583a0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[30]));
  AL_DFF_X al_b3b8ce29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[31]));
  AL_DFF_X al_47d7488b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[32]));
  AL_DFF_X al_25adc2f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[33]));
  AL_DFF_X al_b48349b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[34]));
  AL_DFF_X al_f1df7ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[35]));
  AL_DFF_X al_f858caca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[36]));
  AL_DFF_X al_3452c678 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[37]));
  AL_DFF_X al_15ccfec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[38]));
  AL_DFF_X al_e05382ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[39]));
  AL_DFF_X al_ccb50cd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[40]));
  AL_DFF_X al_c614f60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[41]));
  AL_DFF_X al_a8a86963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[42]));
  AL_DFF_X al_9f4340ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[43]));
  AL_DFF_X al_2cbecf99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[44]));
  AL_DFF_X al_b9dac1b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[45]));
  AL_DFF_X al_dce6434b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[46]));
  AL_DFF_X al_32a5025d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[47]));
  AL_DFF_X al_d5bc18b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[48]));
  AL_DFF_X al_1863740 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[49]));
  AL_DFF_X al_3571e8ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[50]));
  AL_DFF_X al_a613ef49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[51]));
  AL_DFF_X al_f29ed0b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[8]));
  AL_DFF_X al_cd771ed8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[9]));
  AL_DFF_X al_604330b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[10]));
  AL_DFF_X al_3bd284a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[11]));
  AL_DFF_X al_b666db1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[12]));
  AL_DFF_X al_593dd5db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[13]));
  AL_DFF_X al_66c9304f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[14]));
  AL_DFF_X al_6f0de5d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[15]));
  AL_DFF_X al_9b2782fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[16]));
  AL_DFF_X al_ddd48961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[17]));
  AL_DFF_X al_14954d52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[0]));
  AL_DFF_X al_f6c92618 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[18]));
  AL_DFF_X al_26a280a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[19]));
  AL_DFF_X al_d4f76446 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[20]));
  AL_DFF_X al_7ef88d68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[21]));
  AL_DFF_X al_c47faccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[22]));
  AL_DFF_X al_9ae2f727 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[23]));
  AL_DFF_X al_fe0768cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[24]));
  AL_DFF_X al_1d443c73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[25]));
  AL_DFF_X al_e6565a67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[26]));
  AL_DFF_X al_c5abe036 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[27]));
  AL_DFF_X al_418751ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[1]));
  AL_DFF_X al_f1c8e313 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[28]));
  AL_DFF_X al_74e629b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[29]));
  AL_DFF_X al_8058bf2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[30]));
  AL_DFF_X al_9d7a55d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[31]));
  AL_DFF_X al_9dcc0252 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[2]));
  AL_DFF_X al_d85d9278 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[3]));
  AL_DFF_X al_b1620d1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[4]));
  AL_DFF_X al_fcb660bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[5]));
  AL_DFF_X al_c0605feb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[6]));
  AL_DFF_X al_5ea340e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[7]));
  AL_DFF_X al_5f22dd03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[8]));
  AL_DFF_X al_b9009877 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[9]));
  AL_DFF_X al_1b89e8db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[10]));
  AL_DFF_X al_70c9fd7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e3a4cb77),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[0]));
  AL_DFF_X al_83ceed4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[1]));
  AL_DFF_X al_a3c2311e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[2]));
  AL_DFF_X al_b36882d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[3]));
  AL_DFF_X al_b06564c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[4]));
  AL_DFF_X al_ae46ab7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[5]));
  AL_DFF_X al_2da1b0fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[6]));
  AL_DFF_X al_12d06d40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_eac21b5a (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .o(al_42e0e24e));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_7a13e77f (
    .a(1'b0),
    .o({al_6c8e3937,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_895c932f (
    .a(al_6c6869d7[20]),
    .b(al_177a13cd[20]),
    .c(al_6c8e3937),
    .o({al_dbc3e2b0,al_e45a58d8[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5262b9ae (
    .a(al_6c6869d7[21]),
    .b(al_177a13cd[21]),
    .c(al_dbc3e2b0),
    .o({al_a04b98a0,al_e45a58d8[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88524766 (
    .a(al_6c6869d7[22]),
    .b(al_177a13cd[22]),
    .c(al_a04b98a0),
    .o({al_e0aedfd3,al_e45a58d8[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cac3f08 (
    .a(al_6c6869d7[23]),
    .b(al_177a13cd[23]),
    .c(al_e0aedfd3),
    .o({al_150d105b,al_e45a58d8[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_665acdf0 (
    .a(al_6c6869d7[24]),
    .b(al_177a13cd[24]),
    .c(al_150d105b),
    .o({al_6f78cae7,al_e45a58d8[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bdf206d8 (
    .a(al_6c6869d7[25]),
    .b(al_177a13cd[25]),
    .c(al_6f78cae7),
    .o({al_2e62154a,al_e45a58d8[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_65ebca41 (
    .a(al_6c6869d7[26]),
    .b(al_177a13cd[26]),
    .c(al_2e62154a),
    .o({al_e5b9a180,al_e45a58d8[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5206a08 (
    .a(al_6c6869d7[27]),
    .b(al_177a13cd[27]),
    .c(al_e5b9a180),
    .o({al_a4e131c6,al_e45a58d8[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_69065452 (
    .a(al_6c6869d7[28]),
    .b(al_177a13cd[28]),
    .c(al_a4e131c6),
    .o({al_7087d50d,al_e45a58d8[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dba1ec7 (
    .a(al_6c6869d7[29]),
    .b(al_177a13cd[29]),
    .c(al_7087d50d),
    .o({al_6b08641e,al_e45a58d8[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d86e8ba4 (
    .a(al_6c6869d7[30]),
    .b(al_177a13cd[30]),
    .c(al_6b08641e),
    .o({al_b95fb7ea,al_e45a58d8[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92a17348 (
    .a(al_6c6869d7[31]),
    .b(al_177a13cd[31]),
    .c(al_b95fb7ea),
    .o({al_ac18f4f8,al_e45a58d8[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5293decd (
    .c(al_ac18f4f8),
    .o({open_n11,al_e45a58d8[12]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_11887324 (
    .a(al_177a13cd[40]),
    .b(al_177a13cd[41]),
    .c(al_177a13cd[42]),
    .d(al_177a13cd[43]),
    .e(al_177a13cd[44]),
    .f(al_177a13cd[45]),
    .o(al_8cbaef5d));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_5dde944 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[20]),
    .e(al_e45a58d8[0]),
    .o(al_c2901510[20]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_e5bad527 (
    .a(al_177a13cd[48]),
    .b(al_177a13cd[49]),
    .c(al_177a13cd[50]),
    .d(al_177a13cd[51]),
    .o(al_8c892fd7));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_49ed99e (
    .a(al_8cbaef5d),
    .b(al_8c892fd7),
    .c(al_177a13cd[46]),
    .d(al_177a13cd[47]),
    .o(al_eb1649fe));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_af1b52ac (
    .a(al_177a13cd[34]),
    .b(al_177a13cd[35]),
    .c(al_177a13cd[36]),
    .d(al_177a13cd[37]),
    .e(al_177a13cd[38]),
    .f(al_177a13cd[39]),
    .o(al_7b45fe04));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_24c7759b (
    .a(al_177a13cd[32]),
    .b(al_177a13cd[33]),
    .c(al_e45a58d8[12]),
    .o(al_8035eade));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_fe908ac4 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[21]),
    .e(al_e45a58d8[1]),
    .o(al_c2901510[21]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_64e12b76 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[22]),
    .e(al_e45a58d8[2]),
    .o(al_c2901510[22]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_4d98bf1f (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[23]),
    .e(al_e45a58d8[3]),
    .o(al_c2901510[23]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_34f223a4 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[24]),
    .e(al_e45a58d8[4]),
    .o(al_c2901510[24]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_f72e1048 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[25]),
    .e(al_e45a58d8[5]),
    .o(al_c2901510[25]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_2f74844 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[26]),
    .e(al_e45a58d8[6]),
    .o(al_c2901510[26]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_426ebb08 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[27]),
    .e(al_e45a58d8[7]),
    .o(al_c2901510[27]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_cabb262b (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[28]),
    .e(al_e45a58d8[8]),
    .o(al_c2901510[28]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_c662e2ca (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[29]),
    .e(al_e45a58d8[9]),
    .o(al_c2901510[29]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_597ea2be (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[30]),
    .e(al_e45a58d8[10]),
    .o(al_c2901510[30]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_9e50d3c3 (
    .a(al_eb1649fe),
    .b(al_7b45fe04),
    .c(al_8035eade),
    .d(al_6c6869d7[31]),
    .e(al_e45a58d8[11]),
    .o(al_c2901510[31]));
  AL_DFF_X al_5f791956 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_adb04807[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e1bd9dc[0]));
  AL_DFF_X al_34c200c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[19]));
  AL_DFF_X al_bd2400d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[20]));
  AL_DFF_X al_f6697d88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[21]));
  AL_DFF_X al_a32ec72d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[22]));
  AL_DFF_X al_2f9009d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[23]));
  AL_DFF_X al_db253998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[24]));
  AL_DFF_X al_e97b611f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[25]));
  AL_DFF_X al_73b61fe4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[26]));
  AL_DFF_X al_fb929505 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[27]));
  AL_DFF_X al_543ea90c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[28]));
  AL_DFF_X al_d06e794a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[29]));
  AL_DFF_X al_5d9b7d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[30]));
  AL_DFF_X al_8e6ed4cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[31]));
  AL_DFF_X al_526258ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[32]));
  AL_DFF_X al_d0ab0ccc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[33]));
  AL_DFF_X al_1ffb6f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[34]));
  AL_DFF_X al_535bd3b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[35]));
  AL_DFF_X al_fa75ef2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[36]));
  AL_DFF_X al_60fc7e1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[37]));
  AL_DFF_X al_7eea69c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[38]));
  AL_DFF_X al_18e23d10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[39]));
  AL_DFF_X al_ee970a2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[40]));
  AL_DFF_X al_faf51371 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[41]));
  AL_DFF_X al_9fe9a2ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[42]));
  AL_DFF_X al_41f43a98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[43]));
  AL_DFF_X al_e642c1a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[44]));
  AL_DFF_X al_ed7ba649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[45]));
  AL_DFF_X al_83586d3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[46]));
  AL_DFF_X al_fd61660c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[47]));
  AL_DFF_X al_c86c474 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[48]));
  AL_DFF_X al_c33e78e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[49]));
  AL_DFF_X al_ec86df0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[50]));
  AL_DFF_X al_4cf61901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[8]));
  AL_DFF_X al_eed722c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[9]));
  AL_DFF_X al_c103c36f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[10]));
  AL_DFF_X al_304a092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[11]));
  AL_DFF_X al_5af159d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[12]));
  AL_DFF_X al_52ab19ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[13]));
  AL_DFF_X al_d157523b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[14]));
  AL_DFF_X al_c35a923f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[15]));
  AL_DFF_X al_14345ba2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[16]));
  AL_DFF_X al_3f055f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[17]));
  AL_DFF_X al_33dc4ee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[0]));
  AL_DFF_X al_1a3ce8ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[18]));
  AL_DFF_X al_fd8edae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[19]));
  AL_DFF_X al_7fd0e451 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[20]));
  AL_DFF_X al_80037936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[21]));
  AL_DFF_X al_8c913d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[22]));
  AL_DFF_X al_3310d3bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[23]));
  AL_DFF_X al_c84c16e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[24]));
  AL_DFF_X al_7e4881f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[25]));
  AL_DFF_X al_42a3d644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[26]));
  AL_DFF_X al_a4575184 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[27]));
  AL_DFF_X al_fd1a9ca6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[1]));
  AL_DFF_X al_ca7a9ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[28]));
  AL_DFF_X al_52674c79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[29]));
  AL_DFF_X al_35e8fe55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[30]));
  AL_DFF_X al_8d8ff626 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[31]));
  AL_DFF_X al_5f6c3131 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[2]));
  AL_DFF_X al_e3e29066 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[3]));
  AL_DFF_X al_901f2fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[4]));
  AL_DFF_X al_fab4de6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[5]));
  AL_DFF_X al_f080bb8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[6]));
  AL_DFF_X al_e41409eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[7]));
  AL_DFF_X al_9c05d46f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[8]));
  AL_DFF_X al_770bbe03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[9]));
  AL_DFF_X al_2a33c076 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[10]));
  AL_DFF_X al_d0410960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[11]));
  AL_DFF_X al_fc700351 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_42e0e24e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[0]));
  AL_DFF_X al_915e10a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[1]));
  AL_DFF_X al_e76937d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[2]));
  AL_DFF_X al_2ffe15d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[3]));
  AL_DFF_X al_f8dbe566 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[4]));
  AL_DFF_X al_dafcd5c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[5]));
  AL_DFF_X al_7c731645 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[6]));
  AL_DFF_X al_f311d2ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_844d8031 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .o(al_d72d321f));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d4041894 (
    .a(1'b0),
    .o({al_71245cc2,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5bb8a3f (
    .a(al_13d2e70f[19]),
    .b(al_a6f4a789[19]),
    .c(al_71245cc2),
    .o({al_32780627,al_39a3b856[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a2a622d7 (
    .a(al_13d2e70f[20]),
    .b(al_a6f4a789[20]),
    .c(al_32780627),
    .o({al_65eed942,al_39a3b856[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a8eae207 (
    .a(al_13d2e70f[21]),
    .b(al_a6f4a789[21]),
    .c(al_65eed942),
    .o({al_74dcac58,al_39a3b856[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2fbfcb2 (
    .a(al_13d2e70f[22]),
    .b(al_a6f4a789[22]),
    .c(al_74dcac58),
    .o({al_5da4a00d,al_39a3b856[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_df50b67e (
    .a(al_13d2e70f[23]),
    .b(al_a6f4a789[23]),
    .c(al_5da4a00d),
    .o({al_beb32d78,al_39a3b856[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f9b40b3 (
    .a(al_13d2e70f[24]),
    .b(al_a6f4a789[24]),
    .c(al_beb32d78),
    .o({al_32d68c1d,al_39a3b856[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b49d3ec6 (
    .a(al_13d2e70f[25]),
    .b(al_a6f4a789[25]),
    .c(al_32d68c1d),
    .o({al_41f22393,al_39a3b856[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2875dafe (
    .a(al_13d2e70f[26]),
    .b(al_a6f4a789[26]),
    .c(al_41f22393),
    .o({al_28817105,al_39a3b856[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5645f2eb (
    .a(al_13d2e70f[27]),
    .b(al_a6f4a789[27]),
    .c(al_28817105),
    .o({al_93c58a47,al_39a3b856[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fbdb00dd (
    .a(al_13d2e70f[28]),
    .b(al_a6f4a789[28]),
    .c(al_93c58a47),
    .o({al_8b10921e,al_39a3b856[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4baee736 (
    .a(al_13d2e70f[29]),
    .b(al_a6f4a789[29]),
    .c(al_8b10921e),
    .o({al_806ca727,al_39a3b856[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d822766b (
    .a(al_13d2e70f[30]),
    .b(al_a6f4a789[30]),
    .c(al_806ca727),
    .o({al_f4ebe63d,al_39a3b856[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45dc26db (
    .a(al_13d2e70f[31]),
    .b(al_a6f4a789[31]),
    .c(al_f4ebe63d),
    .o({al_b1ae99ca,al_39a3b856[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54f3f6e5 (
    .c(al_b1ae99ca),
    .o({open_n17,al_39a3b856[13]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_22462930 (
    .a(al_a6f4a789[34]),
    .b(al_a6f4a789[35]),
    .c(al_a6f4a789[36]),
    .d(al_a6f4a789[37]),
    .e(al_a6f4a789[38]),
    .f(al_a6f4a789[39]),
    .o(al_c7b36065));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_5fa08e39 (
    .a(al_a6f4a789[42]),
    .b(al_a6f4a789[43]),
    .c(al_a6f4a789[44]),
    .d(al_a6f4a789[45]),
    .o(al_466d66e9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_d4e7d1da (
    .a(al_c7b36065),
    .b(al_466d66e9),
    .c(al_a6f4a789[40]),
    .d(al_a6f4a789[41]),
    .o(al_cb6f9733));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_28f6a66d (
    .a(al_a6f4a789[46]),
    .b(al_a6f4a789[47]),
    .c(al_a6f4a789[48]),
    .d(al_a6f4a789[49]),
    .e(al_a6f4a789[50]),
    .f(al_39a3b856[13]),
    .o(al_884856d));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_7308690c (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[19]),
    .f(al_39a3b856[0]),
    .o(al_fb9cdc0e[19]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_87bab4a6 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[20]),
    .f(al_39a3b856[1]),
    .o(al_fb9cdc0e[20]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_a28b3d1c (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[21]),
    .f(al_39a3b856[2]),
    .o(al_fb9cdc0e[21]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_e58207a9 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[22]),
    .f(al_39a3b856[3]),
    .o(al_fb9cdc0e[22]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_2c33e3b9 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[23]),
    .f(al_39a3b856[4]),
    .o(al_fb9cdc0e[23]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_d93c8308 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[24]),
    .f(al_39a3b856[5]),
    .o(al_fb9cdc0e[24]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_7d77bffc (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[25]),
    .f(al_39a3b856[6]),
    .o(al_fb9cdc0e[25]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_1f0826e5 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[26]),
    .f(al_39a3b856[7]),
    .o(al_fb9cdc0e[26]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_8f706aa1 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[27]),
    .f(al_39a3b856[8]),
    .o(al_fb9cdc0e[27]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_65b22963 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[28]),
    .f(al_39a3b856[9]),
    .o(al_fb9cdc0e[28]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_d8872e4b (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[29]),
    .f(al_39a3b856[10]),
    .o(al_fb9cdc0e[29]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_8e40d222 (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[30]),
    .f(al_39a3b856[11]),
    .o(al_fb9cdc0e[30]));
  AL_MAP_LUT6 #(
    .EQN("(E*~(F)*~((~D*~C*B*A))+E*F*~((~D*~C*B*A))+~(E)*F*(~D*~C*B*A)+E*F*(~D*~C*B*A))"),
    .INIT(64'hffff0008fff70000))
    al_e730aec (
    .a(al_cb6f9733),
    .b(al_884856d),
    .c(al_a6f4a789[32]),
    .d(al_a6f4a789[33]),
    .e(al_13d2e70f[31]),
    .f(al_39a3b856[12]),
    .o(al_fb9cdc0e[31]));
  AL_DFF_X al_aaa8ca34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e1bd9dc[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6d10c98[0]));
  AL_DFF_X al_748f363d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[18]));
  AL_DFF_X al_50f586ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[19]));
  AL_DFF_X al_a23c717a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[20]));
  AL_DFF_X al_ad0a7b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[21]));
  AL_DFF_X al_f5ab502d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[22]));
  AL_DFF_X al_ed7988bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[23]));
  AL_DFF_X al_6f0ab37f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[24]));
  AL_DFF_X al_8dcd789 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[25]));
  AL_DFF_X al_afae7fbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[26]));
  AL_DFF_X al_ee465d46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[27]));
  AL_DFF_X al_6248e6ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[28]));
  AL_DFF_X al_977731c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[29]));
  AL_DFF_X al_aea65d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[30]));
  AL_DFF_X al_ce591abb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[31]));
  AL_DFF_X al_3067931b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[32]));
  AL_DFF_X al_be64ca98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[33]));
  AL_DFF_X al_da4d49f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[34]));
  AL_DFF_X al_7055311f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[35]));
  AL_DFF_X al_88363346 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[36]));
  AL_DFF_X al_9406fa22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[37]));
  AL_DFF_X al_9d11602a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[38]));
  AL_DFF_X al_b6bda817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[39]));
  AL_DFF_X al_abcf3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[40]));
  AL_DFF_X al_84932576 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[41]));
  AL_DFF_X al_1e6f035f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[42]));
  AL_DFF_X al_59312ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[43]));
  AL_DFF_X al_7783c092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[44]));
  AL_DFF_X al_925651f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[45]));
  AL_DFF_X al_c2565f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[46]));
  AL_DFF_X al_c0b11ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[47]));
  AL_DFF_X al_fba6c73d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[48]));
  AL_DFF_X al_d8d7d150 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[49]));
  AL_DFF_X al_2b83ba24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[8]));
  AL_DFF_X al_77f16e1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[9]));
  AL_DFF_X al_fa7cd85e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[10]));
  AL_DFF_X al_a78debcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[11]));
  AL_DFF_X al_c85c958a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[12]));
  AL_DFF_X al_4f71a056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[13]));
  AL_DFF_X al_f7c3a2fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[14]));
  AL_DFF_X al_cb8ed1f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[15]));
  AL_DFF_X al_8e51365d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[16]));
  AL_DFF_X al_faf23c39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[17]));
  AL_DFF_X al_5c601106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[0]));
  AL_DFF_X al_482cf114 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[18]));
  AL_DFF_X al_fd46d3ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[19]));
  AL_DFF_X al_a95b2dca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[20]));
  AL_DFF_X al_c0a7b4d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[21]));
  AL_DFF_X al_225bfd41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[22]));
  AL_DFF_X al_45e5a007 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[23]));
  AL_DFF_X al_b045ce5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[24]));
  AL_DFF_X al_b89b619a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[25]));
  AL_DFF_X al_8356c8ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[26]));
  AL_DFF_X al_1b57e330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[27]));
  AL_DFF_X al_afae26d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[1]));
  AL_DFF_X al_12ccd7cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[28]));
  AL_DFF_X al_78b80428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[29]));
  AL_DFF_X al_e2616c4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[30]));
  AL_DFF_X al_23d7199a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[31]));
  AL_DFF_X al_6a189c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[2]));
  AL_DFF_X al_8053305b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[3]));
  AL_DFF_X al_60e6866b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[4]));
  AL_DFF_X al_e211d44f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[5]));
  AL_DFF_X al_c50f750a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[6]));
  AL_DFF_X al_d43426b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[7]));
  AL_DFF_X al_99372ada (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[8]));
  AL_DFF_X al_bdadbd3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[9]));
  AL_DFF_X al_a5518ac0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[10]));
  AL_DFF_X al_e78a7286 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[11]));
  AL_DFF_X al_819471c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[12]));
  AL_DFF_X al_553eb0e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d72d321f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[0]));
  AL_DFF_X al_b85f7151 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[1]));
  AL_DFF_X al_32b7ffea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[2]));
  AL_DFF_X al_edb277fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[3]));
  AL_DFF_X al_aee99024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[4]));
  AL_DFF_X al_3b900ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[5]));
  AL_DFF_X al_e2c1d6e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[6]));
  AL_DFF_X al_d7e63ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_e26e33bb (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_5ced65c5[14]),
    .o(al_1f755058));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_b31d1d8c (
    .a(1'b0),
    .o({al_5742b37b,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2e4f36a (
    .a(al_7cada4c1[18]),
    .b(al_515b933[18]),
    .c(al_5742b37b),
    .o({al_e4c6cc49,al_5ced65c5[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1a061ada (
    .a(al_7cada4c1[19]),
    .b(al_515b933[19]),
    .c(al_e4c6cc49),
    .o({al_6f18daeb,al_5ced65c5[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8abfe13 (
    .a(al_7cada4c1[20]),
    .b(al_515b933[20]),
    .c(al_6f18daeb),
    .o({al_3fd86060,al_5ced65c5[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7ce51378 (
    .a(al_7cada4c1[21]),
    .b(al_515b933[21]),
    .c(al_3fd86060),
    .o({al_7fd69b02,al_5ced65c5[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e73aab64 (
    .a(al_7cada4c1[22]),
    .b(al_515b933[22]),
    .c(al_7fd69b02),
    .o({al_3b5f5572,al_5ced65c5[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fe94a29 (
    .a(al_7cada4c1[23]),
    .b(al_515b933[23]),
    .c(al_3b5f5572),
    .o({al_926f19c9,al_5ced65c5[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_508c91f2 (
    .a(al_7cada4c1[24]),
    .b(al_515b933[24]),
    .c(al_926f19c9),
    .o({al_71819c0f,al_5ced65c5[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_44ffa8b (
    .a(al_7cada4c1[25]),
    .b(al_515b933[25]),
    .c(al_71819c0f),
    .o({al_16cd5903,al_5ced65c5[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36e91804 (
    .a(al_7cada4c1[26]),
    .b(al_515b933[26]),
    .c(al_16cd5903),
    .o({al_f4b0959f,al_5ced65c5[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b7dedb6 (
    .a(al_7cada4c1[27]),
    .b(al_515b933[27]),
    .c(al_f4b0959f),
    .o({al_b87d9ba8,al_5ced65c5[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f22e747 (
    .a(al_7cada4c1[28]),
    .b(al_515b933[28]),
    .c(al_b87d9ba8),
    .o({al_415da9aa,al_5ced65c5[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f71cfb59 (
    .a(al_7cada4c1[29]),
    .b(al_515b933[29]),
    .c(al_415da9aa),
    .o({al_8465c727,al_5ced65c5[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_965b7e1b (
    .a(al_7cada4c1[30]),
    .b(al_515b933[30]),
    .c(al_8465c727),
    .o({al_f7c19df7,al_5ced65c5[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3042211 (
    .a(al_7cada4c1[31]),
    .b(al_515b933[31]),
    .c(al_f7c19df7),
    .o({al_3ed120c9,al_5ced65c5[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_244f8c2b (
    .c(al_3ed120c9),
    .o({open_n23,al_5ced65c5[14]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_61695e13 (
    .a(al_515b933[38]),
    .b(al_515b933[39]),
    .c(al_515b933[40]),
    .d(al_515b933[41]),
    .e(al_515b933[42]),
    .f(al_515b933[43]),
    .o(al_3f4489bf));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_ef2b84a6 (
    .a(al_515b933[46]),
    .b(al_515b933[47]),
    .c(al_515b933[48]),
    .d(al_515b933[49]),
    .o(al_ae5b1fc6));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_84cadcb9 (
    .a(al_3f4489bf),
    .b(al_ae5b1fc6),
    .c(al_515b933[44]),
    .d(al_515b933[45]),
    .o(al_858ee963));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_71afe415 (
    .a(al_515b933[32]),
    .b(al_515b933[33]),
    .c(al_515b933[34]),
    .d(al_515b933[35]),
    .e(al_515b933[36]),
    .f(al_515b933[37]),
    .o(al_c2097ceb));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_46259cfc (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[18]),
    .d(al_5ced65c5[0]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[18]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_50464ad2 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[19]),
    .d(al_5ced65c5[1]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[19]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_d259c2de (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[20]),
    .d(al_5ced65c5[2]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[20]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_1bfb4587 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[21]),
    .d(al_5ced65c5[3]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[21]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_6b7b00a6 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[22]),
    .d(al_5ced65c5[4]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[22]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_c095dfe7 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[23]),
    .d(al_5ced65c5[5]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[23]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_fc6d485c (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[24]),
    .d(al_5ced65c5[6]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[24]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_bf8fe92d (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[25]),
    .d(al_5ced65c5[7]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[25]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_6dc8104f (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[26]),
    .d(al_5ced65c5[8]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[26]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_b9a2c7d0 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[27]),
    .d(al_5ced65c5[9]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[27]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_41591ed9 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[28]),
    .d(al_5ced65c5[10]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[28]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_4646cd8f (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[29]),
    .d(al_5ced65c5[11]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[29]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_26603a0c (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[30]),
    .d(al_5ced65c5[12]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[30]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D)*~((~E*B*A))+C*D*~((~E*B*A))+~(C)*D*(~E*B*A)+C*D*(~E*B*A))"),
    .INIT(32'hf0f0f870))
    al_e996f628 (
    .a(al_858ee963),
    .b(al_c2097ceb),
    .c(al_7cada4c1[31]),
    .d(al_5ced65c5[13]),
    .e(al_5ced65c5[14]),
    .o(al_28d525d8[31]));
  AL_DFF_X al_f8830cb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c6d10c98[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_599810dd[0]));
  AL_DFF_X al_698ce9b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[17]));
  AL_DFF_X al_fb80e4a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[18]));
  AL_DFF_X al_1c32db03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[19]));
  AL_DFF_X al_b73d4bf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[20]));
  AL_DFF_X al_3728a09b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[21]));
  AL_DFF_X al_bf582eb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[22]));
  AL_DFF_X al_fe1be736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[23]));
  AL_DFF_X al_35a28fa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[24]));
  AL_DFF_X al_76667db4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[25]));
  AL_DFF_X al_e6f03079 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[26]));
  AL_DFF_X al_90ded8ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[27]));
  AL_DFF_X al_5b43e835 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[28]));
  AL_DFF_X al_b60da357 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[29]));
  AL_DFF_X al_c947844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[30]));
  AL_DFF_X al_1bea2287 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[31]));
  AL_DFF_X al_e5503116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[32]));
  AL_DFF_X al_cb7a7dfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[33]));
  AL_DFF_X al_47ae03f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[34]));
  AL_DFF_X al_b44f00c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[35]));
  AL_DFF_X al_431c8d89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[36]));
  AL_DFF_X al_db3a9c3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[37]));
  AL_DFF_X al_b75a9fe4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[38]));
  AL_DFF_X al_dd96ff21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[39]));
  AL_DFF_X al_bfae0d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[40]));
  AL_DFF_X al_38a8598b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[41]));
  AL_DFF_X al_75375c97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[42]));
  AL_DFF_X al_e702ac84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[43]));
  AL_DFF_X al_ea591fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[44]));
  AL_DFF_X al_cb09bb66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[45]));
  AL_DFF_X al_1c3d21af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[46]));
  AL_DFF_X al_e645636f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[47]));
  AL_DFF_X al_50725f0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[48]));
  AL_DFF_X al_86046ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[8]));
  AL_DFF_X al_e557f481 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[9]));
  AL_DFF_X al_b7a0079b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[10]));
  AL_DFF_X al_685631a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[11]));
  AL_DFF_X al_ebbd4b5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[12]));
  AL_DFF_X al_7e56a905 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[13]));
  AL_DFF_X al_323e12f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[14]));
  AL_DFF_X al_f7992c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[15]));
  AL_DFF_X al_5ad021a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[16]));
  AL_DFF_X al_9e431c57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[17]));
  AL_DFF_X al_bdc43bed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[0]));
  AL_DFF_X al_21af9ede (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[18]));
  AL_DFF_X al_64e164ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[19]));
  AL_DFF_X al_16ce962e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[20]));
  AL_DFF_X al_f5d1b500 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[21]));
  AL_DFF_X al_58118609 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[22]));
  AL_DFF_X al_de776835 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[23]));
  AL_DFF_X al_2ce61774 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[24]));
  AL_DFF_X al_7959d511 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[25]));
  AL_DFF_X al_8d19ad41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[26]));
  AL_DFF_X al_12e5b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[27]));
  AL_DFF_X al_d6987f2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[1]));
  AL_DFF_X al_33a089c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[28]));
  AL_DFF_X al_1c4401ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[29]));
  AL_DFF_X al_63ec164f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[30]));
  AL_DFF_X al_ef466ba6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[31]));
  AL_DFF_X al_306a6883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[2]));
  AL_DFF_X al_8e061381 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[3]));
  AL_DFF_X al_90011cc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[4]));
  AL_DFF_X al_800619f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[5]));
  AL_DFF_X al_42c726f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[6]));
  AL_DFF_X al_98fed010 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[7]));
  AL_DFF_X al_5d136a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[8]));
  AL_DFF_X al_25872845 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[9]));
  AL_DFF_X al_d77f91b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[10]));
  AL_DFF_X al_e31d4f46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[11]));
  AL_DFF_X al_24b22567 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[12]));
  AL_DFF_X al_43ee8f03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[13]));
  AL_DFF_X al_ed6f1189 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1f755058),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[0]));
  AL_DFF_X al_9af4782 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[1]));
  AL_DFF_X al_974e227a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[2]));
  AL_DFF_X al_7a250627 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[3]));
  AL_DFF_X al_fd2d782d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[4]));
  AL_DFF_X al_62f71813 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[5]));
  AL_DFF_X al_b8c575 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[6]));
  AL_DFF_X al_4923edca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_581d9bc (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .o(al_6222dcd7));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_c356305c (
    .a(1'b0),
    .o({al_1c729801,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e164e73 (
    .a(al_5fd65077[17]),
    .b(al_82ca84f8[17]),
    .c(al_1c729801),
    .o({al_cc2d4a37,al_51f816c9[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af781034 (
    .a(al_5fd65077[18]),
    .b(al_82ca84f8[18]),
    .c(al_cc2d4a37),
    .o({al_171301db,al_51f816c9[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dc96fd4 (
    .a(al_5fd65077[19]),
    .b(al_82ca84f8[19]),
    .c(al_171301db),
    .o({al_b8a0b712,al_51f816c9[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2fd5a9d (
    .a(al_5fd65077[20]),
    .b(al_82ca84f8[20]),
    .c(al_b8a0b712),
    .o({al_5c73d821,al_51f816c9[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_24bba765 (
    .a(al_5fd65077[21]),
    .b(al_82ca84f8[21]),
    .c(al_5c73d821),
    .o({al_6d30b4d3,al_51f816c9[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e1a4ed81 (
    .a(al_5fd65077[22]),
    .b(al_82ca84f8[22]),
    .c(al_6d30b4d3),
    .o({al_c8e591e5,al_51f816c9[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18011cd8 (
    .a(al_5fd65077[23]),
    .b(al_82ca84f8[23]),
    .c(al_c8e591e5),
    .o({al_ba0cc25,al_51f816c9[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebd200fe (
    .a(al_5fd65077[24]),
    .b(al_82ca84f8[24]),
    .c(al_ba0cc25),
    .o({al_3df74a2f,al_51f816c9[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a56b5cc4 (
    .a(al_5fd65077[25]),
    .b(al_82ca84f8[25]),
    .c(al_3df74a2f),
    .o({al_2265cd1e,al_51f816c9[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d901bf90 (
    .a(al_5fd65077[26]),
    .b(al_82ca84f8[26]),
    .c(al_2265cd1e),
    .o({al_eeaf7eee,al_51f816c9[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ac18c81 (
    .a(al_5fd65077[27]),
    .b(al_82ca84f8[27]),
    .c(al_eeaf7eee),
    .o({al_99a412d5,al_51f816c9[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec6e124b (
    .a(al_5fd65077[28]),
    .b(al_82ca84f8[28]),
    .c(al_99a412d5),
    .o({al_6fc7ef08,al_51f816c9[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a3123573 (
    .a(al_5fd65077[29]),
    .b(al_82ca84f8[29]),
    .c(al_6fc7ef08),
    .o({al_60f2f1ac,al_51f816c9[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa1a956d (
    .a(al_5fd65077[30]),
    .b(al_82ca84f8[30]),
    .c(al_60f2f1ac),
    .o({al_fbd5879f,al_51f816c9[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ccab574a (
    .a(al_5fd65077[31]),
    .b(al_82ca84f8[31]),
    .c(al_fbd5879f),
    .o({al_1800fb32,al_51f816c9[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ca0f986f (
    .c(al_1800fb32),
    .o({open_n29,al_51f816c9[15]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_ea795236 (
    .a(al_82ca84f8[32]),
    .b(al_82ca84f8[33]),
    .c(al_82ca84f8[34]),
    .d(al_82ca84f8[35]),
    .e(al_82ca84f8[36]),
    .f(al_82ca84f8[37]),
    .o(al_6bb8dfe8));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6618b921 (
    .a(al_82ca84f8[40]),
    .b(al_82ca84f8[41]),
    .c(al_82ca84f8[42]),
    .d(al_82ca84f8[43]),
    .o(al_a8cd8f3c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_67948e36 (
    .a(al_6bb8dfe8),
    .b(al_a8cd8f3c),
    .c(al_82ca84f8[38]),
    .d(al_82ca84f8[39]),
    .o(al_d4a26700));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d963cdef (
    .a(al_82ca84f8[44]),
    .b(al_82ca84f8[45]),
    .c(al_82ca84f8[46]),
    .d(al_82ca84f8[47]),
    .e(al_82ca84f8[48]),
    .f(al_51f816c9[15]),
    .o(al_632a2e97));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_2b01b7a5 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[17]),
    .d(al_51f816c9[0]),
    .o(al_8d341179[17]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_1cdbea4a (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[18]),
    .d(al_51f816c9[1]),
    .o(al_8d341179[18]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_991aef48 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[19]),
    .d(al_51f816c9[2]),
    .o(al_8d341179[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_a81a1f0b (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[20]),
    .d(al_51f816c9[3]),
    .o(al_8d341179[20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_f09895bf (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[21]),
    .d(al_51f816c9[4]),
    .o(al_8d341179[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_d082bfc7 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[22]),
    .d(al_51f816c9[5]),
    .o(al_8d341179[22]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_59f7d90b (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[23]),
    .d(al_51f816c9[6]),
    .o(al_8d341179[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_137d7dd8 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[24]),
    .d(al_51f816c9[7]),
    .o(al_8d341179[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_1f31622 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[25]),
    .d(al_51f816c9[8]),
    .o(al_8d341179[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_1a52065b (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[26]),
    .d(al_51f816c9[9]),
    .o(al_8d341179[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9f77fe0e (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[27]),
    .d(al_51f816c9[10]),
    .o(al_8d341179[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9b7bc806 (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[28]),
    .d(al_51f816c9[11]),
    .o(al_8d341179[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_d0d6dd6a (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[29]),
    .d(al_51f816c9[12]),
    .o(al_8d341179[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_3bcb3cce (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[30]),
    .d(al_51f816c9[13]),
    .o(al_8d341179[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ff786a8a (
    .a(al_d4a26700),
    .b(al_632a2e97),
    .c(al_5fd65077[31]),
    .d(al_51f816c9[14]),
    .o(al_8d341179[31]));
  AL_DFF_X al_4053f255 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_599810dd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_903e8807[0]));
  AL_DFF_X al_561cfc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[16]));
  AL_DFF_X al_2c7788b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[17]));
  AL_DFF_X al_7590c6d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[18]));
  AL_DFF_X al_4de2c3b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[19]));
  AL_DFF_X al_495c77c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[20]));
  AL_DFF_X al_a2c58de1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[21]));
  AL_DFF_X al_733117c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[22]));
  AL_DFF_X al_88c4bc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[23]));
  AL_DFF_X al_32b18193 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[24]));
  AL_DFF_X al_e1c66fa4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[25]));
  AL_DFF_X al_1c88f529 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[26]));
  AL_DFF_X al_720d79e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[27]));
  AL_DFF_X al_4effc5af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[28]));
  AL_DFF_X al_17bddc57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[29]));
  AL_DFF_X al_7d03f708 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[30]));
  AL_DFF_X al_4f506710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[31]));
  AL_DFF_X al_8486cfa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[32]));
  AL_DFF_X al_61b2c74c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[33]));
  AL_DFF_X al_d04622d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[34]));
  AL_DFF_X al_44ec27de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[35]));
  AL_DFF_X al_231d1169 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[36]));
  AL_DFF_X al_9be577e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[37]));
  AL_DFF_X al_73ee226c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[38]));
  AL_DFF_X al_a845fc64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[39]));
  AL_DFF_X al_df30f270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[40]));
  AL_DFF_X al_47050022 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[41]));
  AL_DFF_X al_e342d45c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[42]));
  AL_DFF_X al_48298302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[43]));
  AL_DFF_X al_5d51f045 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[44]));
  AL_DFF_X al_3d5047a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[45]));
  AL_DFF_X al_27dfeb38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[46]));
  AL_DFF_X al_d3627933 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[47]));
  AL_DFF_X al_9f431268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[8]));
  AL_DFF_X al_8d13b14a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[9]));
  AL_DFF_X al_72fda091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[10]));
  AL_DFF_X al_2509e888 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[11]));
  AL_DFF_X al_ffd7179a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[12]));
  AL_DFF_X al_c646e435 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[13]));
  AL_DFF_X al_715fa628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[14]));
  AL_DFF_X al_db2376cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[15]));
  AL_DFF_X al_c8c9565b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[16]));
  AL_DFF_X al_9960ebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[17]));
  AL_DFF_X al_ac404f09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[0]));
  AL_DFF_X al_cea0ad81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[18]));
  AL_DFF_X al_e4c2bc78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[19]));
  AL_DFF_X al_5e677b3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[20]));
  AL_DFF_X al_e69be806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[21]));
  AL_DFF_X al_d9f9cbe9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[22]));
  AL_DFF_X al_375fd725 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[23]));
  AL_DFF_X al_ffb37d1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[24]));
  AL_DFF_X al_a403de1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[25]));
  AL_DFF_X al_bcdf86bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[26]));
  AL_DFF_X al_2121876b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[27]));
  AL_DFF_X al_720375c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[1]));
  AL_DFF_X al_8243b19e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[28]));
  AL_DFF_X al_801d3c8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[29]));
  AL_DFF_X al_42006d85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[30]));
  AL_DFF_X al_1dc77ab5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[31]));
  AL_DFF_X al_4d97dff5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[2]));
  AL_DFF_X al_6142e897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[3]));
  AL_DFF_X al_49cd93f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[4]));
  AL_DFF_X al_b7228be4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[5]));
  AL_DFF_X al_c0c7c937 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[6]));
  AL_DFF_X al_2ba445bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[7]));
  AL_DFF_X al_a8aac07e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[8]));
  AL_DFF_X al_ebe57c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[9]));
  AL_DFF_X al_ad7f5102 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[10]));
  AL_DFF_X al_91b1c8af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[11]));
  AL_DFF_X al_f9b1ddea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[12]));
  AL_DFF_X al_5f1a5b9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[13]));
  AL_DFF_X al_b2b929a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[14]));
  AL_DFF_X al_618a14dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6222dcd7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[0]));
  AL_DFF_X al_e6496691 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[1]));
  AL_DFF_X al_ff4b8dcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[2]));
  AL_DFF_X al_b0df242c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[3]));
  AL_DFF_X al_356c2c30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[4]));
  AL_DFF_X al_f75d5799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[5]));
  AL_DFF_X al_1e27b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[6]));
  AL_DFF_X al_5702dab4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e2c0f4f4 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .o(al_c3c604b3));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f0f56325 (
    .a(1'b0),
    .o({al_78a5b5c9,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1eb5d2f2 (
    .a(al_174c5039[16]),
    .b(al_297c219f[16]),
    .c(al_78a5b5c9),
    .o({al_9eeae501,al_bcdd8ff0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_83c48786 (
    .a(al_174c5039[17]),
    .b(al_297c219f[17]),
    .c(al_9eeae501),
    .o({al_c05929c6,al_bcdd8ff0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97d68867 (
    .a(al_174c5039[18]),
    .b(al_297c219f[18]),
    .c(al_c05929c6),
    .o({al_b2191d5e,al_bcdd8ff0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_382461f9 (
    .a(al_174c5039[19]),
    .b(al_297c219f[19]),
    .c(al_b2191d5e),
    .o({al_f7339674,al_bcdd8ff0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47c5debe (
    .a(al_174c5039[20]),
    .b(al_297c219f[20]),
    .c(al_f7339674),
    .o({al_6ded130e,al_bcdd8ff0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_56fb7aa9 (
    .a(al_174c5039[21]),
    .b(al_297c219f[21]),
    .c(al_6ded130e),
    .o({al_467f742e,al_bcdd8ff0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a62037ce (
    .a(al_174c5039[22]),
    .b(al_297c219f[22]),
    .c(al_467f742e),
    .o({al_1cf1391b,al_bcdd8ff0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b039652a (
    .a(al_174c5039[23]),
    .b(al_297c219f[23]),
    .c(al_1cf1391b),
    .o({al_d649f6ed,al_bcdd8ff0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c426a849 (
    .a(al_174c5039[24]),
    .b(al_297c219f[24]),
    .c(al_d649f6ed),
    .o({al_d568756b,al_bcdd8ff0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfb23878 (
    .a(al_174c5039[25]),
    .b(al_297c219f[25]),
    .c(al_d568756b),
    .o({al_3f5f9369,al_bcdd8ff0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c4af1c3d (
    .a(al_174c5039[26]),
    .b(al_297c219f[26]),
    .c(al_3f5f9369),
    .o({al_cad8537e,al_bcdd8ff0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5495635d (
    .a(al_174c5039[27]),
    .b(al_297c219f[27]),
    .c(al_cad8537e),
    .o({al_def1a789,al_bcdd8ff0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57382da8 (
    .a(al_174c5039[28]),
    .b(al_297c219f[28]),
    .c(al_def1a789),
    .o({al_e869e5fb,al_bcdd8ff0[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8170bf06 (
    .a(al_174c5039[29]),
    .b(al_297c219f[29]),
    .c(al_e869e5fb),
    .o({al_38880c22,al_bcdd8ff0[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f9e077fe (
    .a(al_174c5039[30]),
    .b(al_297c219f[30]),
    .c(al_38880c22),
    .o({al_74d32fe0,al_bcdd8ff0[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7a66935d (
    .a(al_174c5039[31]),
    .b(al_297c219f[31]),
    .c(al_74d32fe0),
    .o({al_f930adec,al_bcdd8ff0[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e1f8ee8c (
    .c(al_f930adec),
    .o({open_n35,al_bcdd8ff0[16]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_f07df09f (
    .a(al_297c219f[36]),
    .b(al_297c219f[37]),
    .c(al_297c219f[38]),
    .d(al_297c219f[39]),
    .e(al_297c219f[40]),
    .f(al_297c219f[41]),
    .o(al_3cd6c50e));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8e6a095c (
    .a(al_297c219f[44]),
    .b(al_297c219f[45]),
    .c(al_297c219f[46]),
    .d(al_297c219f[47]),
    .o(al_d4f61208));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_bf37d2e3 (
    .a(al_3cd6c50e),
    .b(al_d4f61208),
    .c(al_297c219f[42]),
    .d(al_297c219f[43]),
    .o(al_cc07f579));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_4739dec3 (
    .a(al_297c219f[32]),
    .b(al_297c219f[33]),
    .c(al_297c219f[34]),
    .d(al_297c219f[35]),
    .e(al_bcdd8ff0[16]),
    .o(al_9d3c2203));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_970ec6ea (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[16]),
    .d(al_bcdd8ff0[0]),
    .o(al_45052583[16]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_aa9bbf44 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[17]),
    .d(al_bcdd8ff0[1]),
    .o(al_45052583[17]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ca13087 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[18]),
    .d(al_bcdd8ff0[2]),
    .o(al_45052583[18]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_f3559c96 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[19]),
    .d(al_bcdd8ff0[3]),
    .o(al_45052583[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_bc13f4b6 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[20]),
    .d(al_bcdd8ff0[4]),
    .o(al_45052583[20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_cf96708b (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[21]),
    .d(al_bcdd8ff0[5]),
    .o(al_45052583[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_a693b417 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[22]),
    .d(al_bcdd8ff0[6]),
    .o(al_45052583[22]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_40bd12e (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[23]),
    .d(al_bcdd8ff0[7]),
    .o(al_45052583[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_94b31228 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[24]),
    .d(al_bcdd8ff0[8]),
    .o(al_45052583[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_317a5d1d (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[25]),
    .d(al_bcdd8ff0[9]),
    .o(al_45052583[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_7a6655a7 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[26]),
    .d(al_bcdd8ff0[10]),
    .o(al_45052583[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9f39cdb8 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[27]),
    .d(al_bcdd8ff0[11]),
    .o(al_45052583[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_fe2f04ec (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[28]),
    .d(al_bcdd8ff0[12]),
    .o(al_45052583[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_22489b67 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[29]),
    .d(al_bcdd8ff0[13]),
    .o(al_45052583[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_6d491d13 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[30]),
    .d(al_bcdd8ff0[14]),
    .o(al_45052583[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_e2753916 (
    .a(al_cc07f579),
    .b(al_9d3c2203),
    .c(al_174c5039[31]),
    .d(al_bcdd8ff0[15]),
    .o(al_45052583[31]));
  AL_DFF_X al_ecd43c29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_903e8807[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5ed5f44b[0]));
  AL_DFF_X al_1d78660c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[15]));
  AL_DFF_X al_46bb5210 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[16]));
  AL_DFF_X al_f762eb32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[17]));
  AL_DFF_X al_1f964a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[18]));
  AL_DFF_X al_d0a6d395 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[19]));
  AL_DFF_X al_5e437793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[20]));
  AL_DFF_X al_473df505 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[21]));
  AL_DFF_X al_adc6e703 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[22]));
  AL_DFF_X al_39faa2c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[23]));
  AL_DFF_X al_30633791 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[24]));
  AL_DFF_X al_6cae4899 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[25]));
  AL_DFF_X al_7032b52b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[26]));
  AL_DFF_X al_28bfd1ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[27]));
  AL_DFF_X al_81853b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[28]));
  AL_DFF_X al_17be0f3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[29]));
  AL_DFF_X al_b4b8e852 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[30]));
  AL_DFF_X al_e1cb120b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[31]));
  AL_DFF_X al_78205801 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[32]));
  AL_DFF_X al_6133919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[33]));
  AL_DFF_X al_ec6b6b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[34]));
  AL_DFF_X al_12439e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[35]));
  AL_DFF_X al_bf4b3d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[36]));
  AL_DFF_X al_cb78feb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[37]));
  AL_DFF_X al_2317e3b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[38]));
  AL_DFF_X al_e55ec464 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[39]));
  AL_DFF_X al_5a4899c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[40]));
  AL_DFF_X al_b8db5cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[41]));
  AL_DFF_X al_efddd755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[42]));
  AL_DFF_X al_96012fb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[43]));
  AL_DFF_X al_670a261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[44]));
  AL_DFF_X al_d61fa757 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[45]));
  AL_DFF_X al_657a10d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[46]));
  AL_DFF_X al_ca7b57a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[8]));
  AL_DFF_X al_69efc6da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[9]));
  AL_DFF_X al_39b51132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[10]));
  AL_DFF_X al_5ad60a25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[11]));
  AL_DFF_X al_4f1ecff0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[12]));
  AL_DFF_X al_8afe9057 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[13]));
  AL_DFF_X al_32d0510d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[14]));
  AL_DFF_X al_9aa3b68f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[15]));
  AL_DFF_X al_3349621b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[16]));
  AL_DFF_X al_bd949bf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[17]));
  AL_DFF_X al_89e7c8ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[0]));
  AL_DFF_X al_346e256c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[18]));
  AL_DFF_X al_871e682b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[19]));
  AL_DFF_X al_d1fd28cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[20]));
  AL_DFF_X al_2b1a37c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[21]));
  AL_DFF_X al_fd0cc140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[22]));
  AL_DFF_X al_d1de55e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[23]));
  AL_DFF_X al_cbb3285c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[24]));
  AL_DFF_X al_27d4a30b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[25]));
  AL_DFF_X al_535f9d7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[26]));
  AL_DFF_X al_606968e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[27]));
  AL_DFF_X al_efd928e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[1]));
  AL_DFF_X al_bc0eaa17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[28]));
  AL_DFF_X al_adf9773d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[29]));
  AL_DFF_X al_ccb8e69d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[30]));
  AL_DFF_X al_b47e36d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[31]));
  AL_DFF_X al_bf5d9e29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[2]));
  AL_DFF_X al_942f8a55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[3]));
  AL_DFF_X al_db5099a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[4]));
  AL_DFF_X al_f3b5ec50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[5]));
  AL_DFF_X al_1a750a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[6]));
  AL_DFF_X al_b8c3846d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[7]));
  AL_DFF_X al_c054bc0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[8]));
  AL_DFF_X al_830ef9ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[9]));
  AL_DFF_X al_353a73a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[10]));
  AL_DFF_X al_676e207c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[11]));
  AL_DFF_X al_4e10cdfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[12]));
  AL_DFF_X al_2261fac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[13]));
  AL_DFF_X al_d452345b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[14]));
  AL_DFF_X al_c90f90ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[15]));
  AL_DFF_X al_fccb916a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c3c604b3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[0]));
  AL_DFF_X al_34f650da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[1]));
  AL_DFF_X al_88474522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[2]));
  AL_DFF_X al_8590dc85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[3]));
  AL_DFF_X al_4fc9bf8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[4]));
  AL_DFF_X al_1378baa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[5]));
  AL_DFF_X al_2876b40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[6]));
  AL_DFF_X al_566840b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_eb7b00ec (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .o(al_5d2d77b4));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_47e1dad4 (
    .a(1'b0),
    .o({al_949714ad,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_199fb287 (
    .a(al_1276f4f7[15]),
    .b(al_2e95330c[15]),
    .c(al_949714ad),
    .o({al_691c6b01,al_d11b8[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_442cf0fc (
    .a(al_1276f4f7[16]),
    .b(al_2e95330c[16]),
    .c(al_691c6b01),
    .o({al_aa40ea6e,al_d11b8[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d196b2ec (
    .a(al_1276f4f7[17]),
    .b(al_2e95330c[17]),
    .c(al_aa40ea6e),
    .o({al_dad76b0c,al_d11b8[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68e10a98 (
    .a(al_1276f4f7[18]),
    .b(al_2e95330c[18]),
    .c(al_dad76b0c),
    .o({al_a0c202f4,al_d11b8[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c5d5eff2 (
    .a(al_1276f4f7[19]),
    .b(al_2e95330c[19]),
    .c(al_a0c202f4),
    .o({al_3ec72efd,al_d11b8[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55fc57e9 (
    .a(al_1276f4f7[20]),
    .b(al_2e95330c[20]),
    .c(al_3ec72efd),
    .o({al_64c5377c,al_d11b8[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a3c12e0 (
    .a(al_1276f4f7[21]),
    .b(al_2e95330c[21]),
    .c(al_64c5377c),
    .o({al_499f819a,al_d11b8[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_134f185e (
    .a(al_1276f4f7[22]),
    .b(al_2e95330c[22]),
    .c(al_499f819a),
    .o({al_d3b6fe74,al_d11b8[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_44b62e8f (
    .a(al_1276f4f7[23]),
    .b(al_2e95330c[23]),
    .c(al_d3b6fe74),
    .o({al_efcf8b1a,al_d11b8[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7db0f264 (
    .a(al_1276f4f7[24]),
    .b(al_2e95330c[24]),
    .c(al_efcf8b1a),
    .o({al_e9939d22,al_d11b8[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3390c684 (
    .a(al_1276f4f7[25]),
    .b(al_2e95330c[25]),
    .c(al_e9939d22),
    .o({al_b2bc9399,al_d11b8[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6e6bb88d (
    .a(al_1276f4f7[26]),
    .b(al_2e95330c[26]),
    .c(al_b2bc9399),
    .o({al_96577a6c,al_d11b8[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae8f3753 (
    .a(al_1276f4f7[27]),
    .b(al_2e95330c[27]),
    .c(al_96577a6c),
    .o({al_a511a420,al_d11b8[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d847c0cf (
    .a(al_1276f4f7[28]),
    .b(al_2e95330c[28]),
    .c(al_a511a420),
    .o({al_523c4f95,al_d11b8[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_301bb555 (
    .a(al_1276f4f7[29]),
    .b(al_2e95330c[29]),
    .c(al_523c4f95),
    .o({al_be2eadc2,al_d11b8[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d23bb395 (
    .a(al_1276f4f7[30]),
    .b(al_2e95330c[30]),
    .c(al_be2eadc2),
    .o({al_1bf3430d,al_d11b8[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_afed7e40 (
    .a(al_1276f4f7[31]),
    .b(al_2e95330c[31]),
    .c(al_1bf3430d),
    .o({al_ee8cd800,al_d11b8[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ea9ca0ac (
    .c(al_ee8cd800),
    .o({open_n41,al_d11b8[17]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_efea26bb (
    .a(al_2e95330c[36]),
    .b(al_2e95330c[37]),
    .c(al_2e95330c[38]),
    .d(al_2e95330c[39]),
    .e(al_2e95330c[40]),
    .f(al_2e95330c[41]),
    .o(al_289b6994));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_4c89ec31 (
    .a(al_2e95330c[44]),
    .b(al_2e95330c[45]),
    .c(al_2e95330c[46]),
    .d(al_d11b8[17]),
    .o(al_278e8e9c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_9bca8c91 (
    .a(al_289b6994),
    .b(al_278e8e9c),
    .c(al_2e95330c[42]),
    .d(al_2e95330c[43]),
    .o(al_62d4794d));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_4bf6136d (
    .a(al_2e95330c[32]),
    .b(al_2e95330c[33]),
    .c(al_2e95330c[34]),
    .d(al_2e95330c[35]),
    .o(al_9d67c14b));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_d02e2ce8 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[15]),
    .d(al_d11b8[0]),
    .o(al_b5df9b8a[15]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_141331c8 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[16]),
    .d(al_d11b8[1]),
    .o(al_b5df9b8a[16]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_17e1b060 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[17]),
    .d(al_d11b8[2]),
    .o(al_b5df9b8a[17]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_555a9a70 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[18]),
    .d(al_d11b8[3]),
    .o(al_b5df9b8a[18]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_42e1ed76 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[19]),
    .d(al_d11b8[4]),
    .o(al_b5df9b8a[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_5e0d4b3c (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[20]),
    .d(al_d11b8[5]),
    .o(al_b5df9b8a[20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_d1f55f22 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[21]),
    .d(al_d11b8[6]),
    .o(al_b5df9b8a[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ab067bbe (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[22]),
    .d(al_d11b8[7]),
    .o(al_b5df9b8a[22]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_5eb34362 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[23]),
    .d(al_d11b8[8]),
    .o(al_b5df9b8a[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_29989d9e (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[24]),
    .d(al_d11b8[9]),
    .o(al_b5df9b8a[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ecc6e306 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[25]),
    .d(al_d11b8[10]),
    .o(al_b5df9b8a[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_15331e5c (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[26]),
    .d(al_d11b8[11]),
    .o(al_b5df9b8a[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_bb16527b (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[27]),
    .d(al_d11b8[12]),
    .o(al_b5df9b8a[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9c44441a (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[28]),
    .d(al_d11b8[13]),
    .o(al_b5df9b8a[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_963f7f04 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[29]),
    .d(al_d11b8[14]),
    .o(al_b5df9b8a[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_11dd5145 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[30]),
    .d(al_d11b8[15]),
    .o(al_b5df9b8a[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_14a69f62 (
    .a(al_62d4794d),
    .b(al_9d67c14b),
    .c(al_1276f4f7[31]),
    .d(al_d11b8[16]),
    .o(al_b5df9b8a[31]));
  AL_DFF_X al_8863fafc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5ed5f44b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_54284e1f[0]));
  AL_DFF_X al_da690016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[14]));
  AL_DFF_X al_2913d12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[15]));
  AL_DFF_X al_f38c9059 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[16]));
  AL_DFF_X al_5c986209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[17]));
  AL_DFF_X al_38c0452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[18]));
  AL_DFF_X al_df3866bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[19]));
  AL_DFF_X al_ece1684 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[20]));
  AL_DFF_X al_dc2f7076 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[21]));
  AL_DFF_X al_3d965b8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[22]));
  AL_DFF_X al_b290a350 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[23]));
  AL_DFF_X al_86a85a01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[24]));
  AL_DFF_X al_e882956e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[25]));
  AL_DFF_X al_7800a95b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[26]));
  AL_DFF_X al_15c5372b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[27]));
  AL_DFF_X al_6bbeef3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[28]));
  AL_DFF_X al_1afe138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[29]));
  AL_DFF_X al_dd24357e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[30]));
  AL_DFF_X al_aacb3bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[31]));
  AL_DFF_X al_cd8faff0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[32]));
  AL_DFF_X al_e4217e2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[33]));
  AL_DFF_X al_f2216d79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[34]));
  AL_DFF_X al_7fd65221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[35]));
  AL_DFF_X al_fa1c10cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[36]));
  AL_DFF_X al_bd389b66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[37]));
  AL_DFF_X al_413a4897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[38]));
  AL_DFF_X al_a8243dec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[39]));
  AL_DFF_X al_c964ab4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[40]));
  AL_DFF_X al_5b7f18e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[41]));
  AL_DFF_X al_bff9eb98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[42]));
  AL_DFF_X al_65c83562 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[43]));
  AL_DFF_X al_218b2cba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[44]));
  AL_DFF_X al_7254a75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[45]));
  AL_DFF_X al_f9204cef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[8]));
  AL_DFF_X al_cdc24628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[9]));
  AL_DFF_X al_e713d18f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[10]));
  AL_DFF_X al_504cc943 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[11]));
  AL_DFF_X al_4f9dbbcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[12]));
  AL_DFF_X al_d74c20e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[13]));
  AL_DFF_X al_445df5ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[14]));
  AL_DFF_X al_cad707e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[15]));
  AL_DFF_X al_e250c528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[16]));
  AL_DFF_X al_d2daa6e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[17]));
  AL_DFF_X al_6648f4e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[0]));
  AL_DFF_X al_c001cb03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[18]));
  AL_DFF_X al_adcc4124 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[19]));
  AL_DFF_X al_eb6298f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[20]));
  AL_DFF_X al_3cacee2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[21]));
  AL_DFF_X al_b69c4a63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[22]));
  AL_DFF_X al_cf5c6ce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[23]));
  AL_DFF_X al_60ead5ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[24]));
  AL_DFF_X al_cdec21fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[25]));
  AL_DFF_X al_a6d08be1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[26]));
  AL_DFF_X al_fc6e3937 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[27]));
  AL_DFF_X al_889833c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[1]));
  AL_DFF_X al_ad2601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[28]));
  AL_DFF_X al_c4cfb66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[29]));
  AL_DFF_X al_ff5872f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[30]));
  AL_DFF_X al_1f74db12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[31]));
  AL_DFF_X al_5db6d60b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[2]));
  AL_DFF_X al_8ab8b26c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[3]));
  AL_DFF_X al_f0ae4188 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[4]));
  AL_DFF_X al_44f5b5e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[5]));
  AL_DFF_X al_fa962868 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[6]));
  AL_DFF_X al_870f6263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[7]));
  AL_DFF_X al_6a3b497b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[8]));
  AL_DFF_X al_bf41ec8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[9]));
  AL_DFF_X al_bfb52963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[10]));
  AL_DFF_X al_be6eb2e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[11]));
  AL_DFF_X al_932ec8c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[12]));
  AL_DFF_X al_e1786ae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[13]));
  AL_DFF_X al_e230a7d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[14]));
  AL_DFF_X al_2d852ba3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[15]));
  AL_DFF_X al_6ac43263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[16]));
  AL_DFF_X al_b035928a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d2d77b4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[0]));
  AL_DFF_X al_8ddaaf4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[1]));
  AL_DFF_X al_658b8325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[2]));
  AL_DFF_X al_4b60cc8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[3]));
  AL_DFF_X al_5fa1ac81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[4]));
  AL_DFF_X al_29653411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[5]));
  AL_DFF_X al_12826897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[6]));
  AL_DFF_X al_8bdc4811 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_e87a18a0 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_2bcf47f2[18]),
    .o(al_579fe9c9));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_e5fe5611 (
    .a(1'b0),
    .o({al_37d85dd8,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_adf63d31 (
    .a(al_3692f86e[14]),
    .b(al_b4e2b23b[14]),
    .c(al_37d85dd8),
    .o({al_22c0f879,al_2bcf47f2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dee5dd53 (
    .a(al_3692f86e[15]),
    .b(al_b4e2b23b[15]),
    .c(al_22c0f879),
    .o({al_a6323dfd,al_2bcf47f2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21726e66 (
    .a(al_3692f86e[16]),
    .b(al_b4e2b23b[16]),
    .c(al_a6323dfd),
    .o({al_d459fd2a,al_2bcf47f2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ed725db (
    .a(al_3692f86e[17]),
    .b(al_b4e2b23b[17]),
    .c(al_d459fd2a),
    .o({al_a0f8478c,al_2bcf47f2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_595cf5e1 (
    .a(al_3692f86e[18]),
    .b(al_b4e2b23b[18]),
    .c(al_a0f8478c),
    .o({al_67dd1cc2,al_2bcf47f2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9f4e33a (
    .a(al_3692f86e[19]),
    .b(al_b4e2b23b[19]),
    .c(al_67dd1cc2),
    .o({al_9380c67b,al_2bcf47f2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fdc966af (
    .a(al_3692f86e[20]),
    .b(al_b4e2b23b[20]),
    .c(al_9380c67b),
    .o({al_6b7d50a7,al_2bcf47f2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a8e8963 (
    .a(al_3692f86e[21]),
    .b(al_b4e2b23b[21]),
    .c(al_6b7d50a7),
    .o({al_4cc7f121,al_2bcf47f2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40fc16b2 (
    .a(al_3692f86e[22]),
    .b(al_b4e2b23b[22]),
    .c(al_4cc7f121),
    .o({al_648c2518,al_2bcf47f2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e250c835 (
    .a(al_3692f86e[23]),
    .b(al_b4e2b23b[23]),
    .c(al_648c2518),
    .o({al_1ba5074a,al_2bcf47f2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b64e2f0e (
    .a(al_3692f86e[24]),
    .b(al_b4e2b23b[24]),
    .c(al_1ba5074a),
    .o({al_959737fa,al_2bcf47f2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_817a3c84 (
    .a(al_3692f86e[25]),
    .b(al_b4e2b23b[25]),
    .c(al_959737fa),
    .o({al_456e9f5b,al_2bcf47f2[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e4ac0b07 (
    .a(al_3692f86e[26]),
    .b(al_b4e2b23b[26]),
    .c(al_456e9f5b),
    .o({al_983289c4,al_2bcf47f2[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_74ef5355 (
    .a(al_3692f86e[27]),
    .b(al_b4e2b23b[27]),
    .c(al_983289c4),
    .o({al_170bfe43,al_2bcf47f2[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fe62cdc2 (
    .a(al_3692f86e[28]),
    .b(al_b4e2b23b[28]),
    .c(al_170bfe43),
    .o({al_96c24183,al_2bcf47f2[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e355d2e6 (
    .a(al_3692f86e[29]),
    .b(al_b4e2b23b[29]),
    .c(al_96c24183),
    .o({al_a7a2d586,al_2bcf47f2[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dc00befa (
    .a(al_3692f86e[30]),
    .b(al_b4e2b23b[30]),
    .c(al_a7a2d586),
    .o({al_1ba7203c,al_2bcf47f2[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_79d4deb2 (
    .a(al_3692f86e[31]),
    .b(al_b4e2b23b[31]),
    .c(al_1ba7203c),
    .o({al_fdbea65d,al_2bcf47f2[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c67fe61d (
    .c(al_fdbea65d),
    .o({open_n47,al_2bcf47f2[18]}));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_df968e04 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[14]),
    .e(al_2bcf47f2[0]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[14]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_73d332c3 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[15]),
    .e(al_2bcf47f2[1]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[15]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d61b036 (
    .a(al_b4e2b23b[34]),
    .b(al_b4e2b23b[35]),
    .c(al_b4e2b23b[36]),
    .d(al_b4e2b23b[37]),
    .e(al_b4e2b23b[38]),
    .f(al_b4e2b23b[39]),
    .o(al_92ca20ed));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d22cc882 (
    .a(al_b4e2b23b[42]),
    .b(al_b4e2b23b[43]),
    .c(al_b4e2b23b[44]),
    .d(al_b4e2b23b[45]),
    .o(al_2758bb5));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_8a6aca2d (
    .a(al_92ca20ed),
    .b(al_2758bb5),
    .c(al_b4e2b23b[40]),
    .d(al_b4e2b23b[41]),
    .o(al_337113ba));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_b6f6ca36 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[16]),
    .e(al_2bcf47f2[2]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[16]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_a464ed60 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[17]),
    .e(al_2bcf47f2[3]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[17]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_8285ca09 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[18]),
    .e(al_2bcf47f2[4]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[18]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_9b6e34e5 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[19]),
    .e(al_2bcf47f2[5]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[19]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_6733f951 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[20]),
    .e(al_2bcf47f2[6]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[20]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_c0f664c9 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[21]),
    .e(al_2bcf47f2[7]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[21]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_69e7dcfc (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[22]),
    .e(al_2bcf47f2[8]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[22]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_9d81a8ca (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[23]),
    .e(al_2bcf47f2[9]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[23]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_636bd497 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[24]),
    .e(al_2bcf47f2[10]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[24]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_628f97b7 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[25]),
    .e(al_2bcf47f2[11]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[25]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_bb4b1448 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[26]),
    .e(al_2bcf47f2[12]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[26]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_b70ef665 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[27]),
    .e(al_2bcf47f2[13]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[27]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_6e31a77b (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[28]),
    .e(al_2bcf47f2[14]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[28]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_e5242341 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[29]),
    .e(al_2bcf47f2[15]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[29]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_85f25e31 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[30]),
    .e(al_2bcf47f2[16]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[30]));
  AL_MAP_LUT6 #(
    .EQN("(D*~(E)*~((~F*~C*~B*A))+D*E*~((~F*~C*~B*A))+~(D)*E*(~F*~C*~B*A)+D*E*(~F*~C*~B*A))"),
    .INIT(64'hff00ff00ff02fd00))
    al_5542f9f5 (
    .a(al_337113ba),
    .b(al_b4e2b23b[32]),
    .c(al_b4e2b23b[33]),
    .d(al_3692f86e[31]),
    .e(al_2bcf47f2[17]),
    .f(al_2bcf47f2[18]),
    .o(al_28955387[31]));
  AL_DFF_X al_c347a0ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_54284e1f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f83a6cd4[0]));
  AL_DFF_X al_1ac62b61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[13]));
  AL_DFF_X al_600f65f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[14]));
  AL_DFF_X al_af6de916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[15]));
  AL_DFF_X al_26879b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[16]));
  AL_DFF_X al_96264659 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[17]));
  AL_DFF_X al_f850b737 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[18]));
  AL_DFF_X al_57025d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[19]));
  AL_DFF_X al_8d2f05eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[20]));
  AL_DFF_X al_86d9eefd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[21]));
  AL_DFF_X al_f4ae2360 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[22]));
  AL_DFF_X al_a7827892 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[23]));
  AL_DFF_X al_da2f76e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[24]));
  AL_DFF_X al_fb5c48fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[25]));
  AL_DFF_X al_e611135d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[26]));
  AL_DFF_X al_dde02ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[27]));
  AL_DFF_X al_fcdddf35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[28]));
  AL_DFF_X al_781abdfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[29]));
  AL_DFF_X al_b2acdef1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[30]));
  AL_DFF_X al_a708b47e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[31]));
  AL_DFF_X al_a76d9052 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[32]));
  AL_DFF_X al_ec26ffc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[33]));
  AL_DFF_X al_10ea39c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[34]));
  AL_DFF_X al_b1215e2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[35]));
  AL_DFF_X al_335e8232 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[36]));
  AL_DFF_X al_e7b392ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[37]));
  AL_DFF_X al_ec02c66b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[38]));
  AL_DFF_X al_c6fb9ac5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[39]));
  AL_DFF_X al_be9d98cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[40]));
  AL_DFF_X al_1393a042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[41]));
  AL_DFF_X al_67b47477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[42]));
  AL_DFF_X al_13dc88ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[43]));
  AL_DFF_X al_6f2d8411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[44]));
  AL_DFF_X al_f282934e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[8]));
  AL_DFF_X al_707b7784 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[9]));
  AL_DFF_X al_598b85d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[10]));
  AL_DFF_X al_8650a834 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[11]));
  AL_DFF_X al_2dab9f6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[12]));
  AL_DFF_X al_8f2ce4ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[13]));
  AL_DFF_X al_f04f456f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[14]));
  AL_DFF_X al_1b064a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[15]));
  AL_DFF_X al_d588437d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[16]));
  AL_DFF_X al_4cb306ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[17]));
  AL_DFF_X al_2c51f322 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[0]));
  AL_DFF_X al_cb30847d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[18]));
  AL_DFF_X al_d861793b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[19]));
  AL_DFF_X al_1573330b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[20]));
  AL_DFF_X al_66a54e9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[21]));
  AL_DFF_X al_bc7e578b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[22]));
  AL_DFF_X al_cae3a25a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[23]));
  AL_DFF_X al_66e905ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[24]));
  AL_DFF_X al_9412a09a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[25]));
  AL_DFF_X al_a81a4530 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[26]));
  AL_DFF_X al_653bc7ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[27]));
  AL_DFF_X al_e9984b4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[1]));
  AL_DFF_X al_49885406 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[28]));
  AL_DFF_X al_3fd661be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[29]));
  AL_DFF_X al_2b901dc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[30]));
  AL_DFF_X al_a4ba2241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[31]));
  AL_DFF_X al_da34ba3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[2]));
  AL_DFF_X al_21e11f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[3]));
  AL_DFF_X al_54732186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[4]));
  AL_DFF_X al_d740ee5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[5]));
  AL_DFF_X al_c724a07b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[6]));
  AL_DFF_X al_5fc5d4a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[7]));
  AL_DFF_X al_40e8250c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[8]));
  AL_DFF_X al_69bc6fa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[9]));
  AL_DFF_X al_32af8f6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[10]));
  AL_DFF_X al_6ee217c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[11]));
  AL_DFF_X al_8d9df29f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[12]));
  AL_DFF_X al_f5433ea7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[13]));
  AL_DFF_X al_b89151a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[14]));
  AL_DFF_X al_55aadca4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[15]));
  AL_DFF_X al_7b5299a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[16]));
  AL_DFF_X al_371816c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[17]));
  AL_DFF_X al_3779d9fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_579fe9c9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[0]));
  AL_DFF_X al_ff1bc292 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[1]));
  AL_DFF_X al_1c758035 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[2]));
  AL_DFF_X al_88819cb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[3]));
  AL_DFF_X al_b48ef4f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[4]));
  AL_DFF_X al_fe001b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[5]));
  AL_DFF_X al_1d7bd91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[6]));
  AL_DFF_X al_34efbac9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_cc8fd5ad (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .o(al_877d1bc));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_c4b9631d (
    .a(1'b0),
    .o({al_b98fe565,open_n50}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86bd31da (
    .a(al_368cfa5b[13]),
    .b(al_e7d838f[13]),
    .c(al_b98fe565),
    .o({al_60ed0a3f,al_f57e3792[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33d49e71 (
    .a(al_368cfa5b[14]),
    .b(al_e7d838f[14]),
    .c(al_60ed0a3f),
    .o({al_27d9400d,al_f57e3792[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_95366194 (
    .a(al_368cfa5b[15]),
    .b(al_e7d838f[15]),
    .c(al_27d9400d),
    .o({al_94badae1,al_f57e3792[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f51c2e7 (
    .a(al_368cfa5b[16]),
    .b(al_e7d838f[16]),
    .c(al_94badae1),
    .o({al_462fcfec,al_f57e3792[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d930076 (
    .a(al_368cfa5b[17]),
    .b(al_e7d838f[17]),
    .c(al_462fcfec),
    .o({al_11444b05,al_f57e3792[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de464f39 (
    .a(al_368cfa5b[18]),
    .b(al_e7d838f[18]),
    .c(al_11444b05),
    .o({al_6a490a84,al_f57e3792[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84d3b065 (
    .a(al_368cfa5b[19]),
    .b(al_e7d838f[19]),
    .c(al_6a490a84),
    .o({al_7c4effa7,al_f57e3792[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_20233178 (
    .a(al_368cfa5b[20]),
    .b(al_e7d838f[20]),
    .c(al_7c4effa7),
    .o({al_2a54b225,al_f57e3792[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_179b2a11 (
    .a(al_368cfa5b[21]),
    .b(al_e7d838f[21]),
    .c(al_2a54b225),
    .o({al_bf2e29ab,al_f57e3792[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_91b4969a (
    .a(al_368cfa5b[22]),
    .b(al_e7d838f[22]),
    .c(al_bf2e29ab),
    .o({al_1741bada,al_f57e3792[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eea1df1d (
    .a(al_368cfa5b[23]),
    .b(al_e7d838f[23]),
    .c(al_1741bada),
    .o({al_506041c3,al_f57e3792[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f4b90e54 (
    .a(al_368cfa5b[24]),
    .b(al_e7d838f[24]),
    .c(al_506041c3),
    .o({al_ff00a5b,al_f57e3792[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a16ded5d (
    .a(al_368cfa5b[25]),
    .b(al_e7d838f[25]),
    .c(al_ff00a5b),
    .o({al_cadab979,al_f57e3792[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_338029f (
    .a(al_368cfa5b[26]),
    .b(al_e7d838f[26]),
    .c(al_cadab979),
    .o({al_1ca453a8,al_f57e3792[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_578a3fe3 (
    .a(al_368cfa5b[27]),
    .b(al_e7d838f[27]),
    .c(al_1ca453a8),
    .o({al_a7dd3d61,al_f57e3792[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a8d670e (
    .a(al_368cfa5b[28]),
    .b(al_e7d838f[28]),
    .c(al_a7dd3d61),
    .o({al_f0c84e95,al_f57e3792[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6bd3f77 (
    .a(al_368cfa5b[29]),
    .b(al_e7d838f[29]),
    .c(al_f0c84e95),
    .o({al_11666a8e,al_f57e3792[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a4c8e1a3 (
    .a(al_368cfa5b[30]),
    .b(al_e7d838f[30]),
    .c(al_11666a8e),
    .o({al_2f88a0b8,al_f57e3792[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_62bc376 (
    .a(al_368cfa5b[31]),
    .b(al_e7d838f[31]),
    .c(al_2f88a0b8),
    .o({al_6a534ff7,al_f57e3792[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_237b3aff (
    .c(al_6a534ff7),
    .o({open_n53,al_f57e3792[19]}));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_3b2d9ee5 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[13]),
    .e(al_f57e3792[0]),
    .o(al_e55e130b[13]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_d7a96bd6 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[14]),
    .e(al_f57e3792[1]),
    .o(al_e55e130b[14]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_cc03f8a7 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[15]),
    .e(al_f57e3792[2]),
    .o(al_e55e130b[15]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_a11bea05 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[16]),
    .e(al_f57e3792[3]),
    .o(al_e55e130b[16]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6bccec7d (
    .a(al_e7d838f[34]),
    .b(al_e7d838f[35]),
    .c(al_e7d838f[36]),
    .d(al_e7d838f[37]),
    .e(al_e7d838f[38]),
    .f(al_e7d838f[39]),
    .o(al_22cba5b6));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_253eb6f (
    .a(al_e7d838f[42]),
    .b(al_e7d838f[43]),
    .c(al_e7d838f[44]),
    .d(al_f57e3792[19]),
    .o(al_dc8a8f4));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_487830fd (
    .a(al_22cba5b6),
    .b(al_dc8a8f4),
    .c(al_e7d838f[40]),
    .d(al_e7d838f[41]),
    .o(al_3ad2f5fe));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_3da221d3 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[17]),
    .e(al_f57e3792[4]),
    .o(al_e55e130b[17]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_b6d26ed3 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[18]),
    .e(al_f57e3792[5]),
    .o(al_e55e130b[18]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_a5bb8a2 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[19]),
    .e(al_f57e3792[6]),
    .o(al_e55e130b[19]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_fdfcb8ec (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[20]),
    .e(al_f57e3792[7]),
    .o(al_e55e130b[20]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_20a0499c (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[21]),
    .e(al_f57e3792[8]),
    .o(al_e55e130b[21]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_a11d1933 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[22]),
    .e(al_f57e3792[9]),
    .o(al_e55e130b[22]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_c4ee51a8 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[23]),
    .e(al_f57e3792[10]),
    .o(al_e55e130b[23]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_9a762858 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[24]),
    .e(al_f57e3792[11]),
    .o(al_e55e130b[24]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_119f1b42 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[25]),
    .e(al_f57e3792[12]),
    .o(al_e55e130b[25]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_e56059a4 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[26]),
    .e(al_f57e3792[13]),
    .o(al_e55e130b[26]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_83588894 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[27]),
    .e(al_f57e3792[14]),
    .o(al_e55e130b[27]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_5ec3ec62 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[28]),
    .e(al_f57e3792[15]),
    .o(al_e55e130b[28]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_b14aa975 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[29]),
    .e(al_f57e3792[16]),
    .o(al_e55e130b[29]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_ee3a7ce4 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[30]),
    .e(al_f57e3792[17]),
    .o(al_e55e130b[30]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~C*~B*A))+D*E*~((~C*~B*A))+~(D)*E*(~C*~B*A)+D*E*(~C*~B*A))"),
    .INIT(32'hff02fd00))
    al_f2b14a41 (
    .a(al_3ad2f5fe),
    .b(al_e7d838f[32]),
    .c(al_e7d838f[33]),
    .d(al_368cfa5b[31]),
    .e(al_f57e3792[18]),
    .o(al_e55e130b[31]));
  AL_DFF_X al_7c9d1b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f83a6cd4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a2efb7[0]));
  AL_DFF_X al_480e70af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[12]));
  AL_DFF_X al_6ce5151d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[13]));
  AL_DFF_X al_275bb04c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[14]));
  AL_DFF_X al_c5a1e024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[15]));
  AL_DFF_X al_5de54e04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[16]));
  AL_DFF_X al_b99a429a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[17]));
  AL_DFF_X al_485e69c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[18]));
  AL_DFF_X al_803d743b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[19]));
  AL_DFF_X al_34a20e08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[20]));
  AL_DFF_X al_4d24a13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[21]));
  AL_DFF_X al_2c3f8dab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[22]));
  AL_DFF_X al_be94bed4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[23]));
  AL_DFF_X al_930dc506 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[24]));
  AL_DFF_X al_f64d2945 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[25]));
  AL_DFF_X al_5ec3c261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[26]));
  AL_DFF_X al_7769fdbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[27]));
  AL_DFF_X al_9b763698 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[28]));
  AL_DFF_X al_55f38d3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[29]));
  AL_DFF_X al_f3edfdb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[30]));
  AL_DFF_X al_59c676e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[31]));
  AL_DFF_X al_b626b137 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[32]));
  AL_DFF_X al_dd4c256c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[33]));
  AL_DFF_X al_9af4d647 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[34]));
  AL_DFF_X al_a600435a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[35]));
  AL_DFF_X al_eaab1171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[36]));
  AL_DFF_X al_a9456a01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[37]));
  AL_DFF_X al_6917ea78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[38]));
  AL_DFF_X al_d141daf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[39]));
  AL_DFF_X al_5742a289 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[40]));
  AL_DFF_X al_d71f8f72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[41]));
  AL_DFF_X al_5bcb02a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[42]));
  AL_DFF_X al_bc0ec360 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[43]));
  AL_DFF_X al_f25143fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[8]));
  AL_DFF_X al_b9a97130 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[9]));
  AL_DFF_X al_59c85dcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[10]));
  AL_DFF_X al_38ceddb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[11]));
  AL_DFF_X al_485caf90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[12]));
  AL_DFF_X al_c12b4419 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[13]));
  AL_DFF_X al_dbdf230c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[14]));
  AL_DFF_X al_d34f3cf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[15]));
  AL_DFF_X al_e674ba6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[16]));
  AL_DFF_X al_99ab243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[17]));
  AL_DFF_X al_769994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[0]));
  AL_DFF_X al_d19d7a8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[18]));
  AL_DFF_X al_460528b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[19]));
  AL_DFF_X al_8b97dcfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[20]));
  AL_DFF_X al_880d91f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[21]));
  AL_DFF_X al_ca650997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[22]));
  AL_DFF_X al_58c93826 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[23]));
  AL_DFF_X al_1c516e37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[24]));
  AL_DFF_X al_ed2820f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[25]));
  AL_DFF_X al_ee428f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[26]));
  AL_DFF_X al_827bf6c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[27]));
  AL_DFF_X al_16ccc308 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[1]));
  AL_DFF_X al_d2889bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[28]));
  AL_DFF_X al_cfbb93a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[29]));
  AL_DFF_X al_e2684f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[30]));
  AL_DFF_X al_5836c2a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[31]));
  AL_DFF_X al_a310666b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[2]));
  AL_DFF_X al_32c6279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[3]));
  AL_DFF_X al_b3908cfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[4]));
  AL_DFF_X al_67adc5ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[5]));
  AL_DFF_X al_f66bd97d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[6]));
  AL_DFF_X al_c25ec0bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[7]));
  AL_DFF_X al_f50ee1eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[8]));
  AL_DFF_X al_4a59c974 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[9]));
  AL_DFF_X al_389be8fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[10]));
  AL_DFF_X al_5b7b006d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[11]));
  AL_DFF_X al_91b528d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[12]));
  AL_DFF_X al_14aa126e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[13]));
  AL_DFF_X al_9353cc3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[14]));
  AL_DFF_X al_2bae2f04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[15]));
  AL_DFF_X al_896875b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[16]));
  AL_DFF_X al_58ad814a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[17]));
  AL_DFF_X al_297837a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_877d1bc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[0]));
  AL_DFF_X al_8611f253 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[18]));
  AL_DFF_X al_d0657014 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[1]));
  AL_DFF_X al_2472a8e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[2]));
  AL_DFF_X al_63765d60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[3]));
  AL_DFF_X al_53ca59e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[4]));
  AL_DFF_X al_602ebf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[5]));
  AL_DFF_X al_49be09d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[6]));
  AL_DFF_X al_5bece1f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_6b118967 (
    .a(al_e8916352),
    .b(al_755dcbd4[20]),
    .o(al_cc19a77c));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1f07a30e (
    .a(1'b0),
    .o({al_80347035,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_61113f9a (
    .a(al_e240f99f[12]),
    .b(al_30e951fe[12]),
    .c(al_80347035),
    .o({al_54975822,al_755dcbd4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e68718e0 (
    .a(al_e240f99f[13]),
    .b(al_30e951fe[13]),
    .c(al_54975822),
    .o({al_e5f75e51,al_755dcbd4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1ffa79 (
    .a(al_e240f99f[14]),
    .b(al_30e951fe[14]),
    .c(al_e5f75e51),
    .o({al_84743aea,al_755dcbd4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b08ab490 (
    .a(al_e240f99f[15]),
    .b(al_30e951fe[15]),
    .c(al_84743aea),
    .o({al_4c6c1136,al_755dcbd4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9ba0fd6c (
    .a(al_e240f99f[16]),
    .b(al_30e951fe[16]),
    .c(al_4c6c1136),
    .o({al_aff6af71,al_755dcbd4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57ba3a96 (
    .a(al_e240f99f[17]),
    .b(al_30e951fe[17]),
    .c(al_aff6af71),
    .o({al_786cd6fa,al_755dcbd4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d29c057c (
    .a(al_e240f99f[18]),
    .b(al_30e951fe[18]),
    .c(al_786cd6fa),
    .o({al_ea94f7fb,al_755dcbd4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fff76b36 (
    .a(al_e240f99f[19]),
    .b(al_30e951fe[19]),
    .c(al_ea94f7fb),
    .o({al_83614d40,al_755dcbd4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_85621d7b (
    .a(al_e240f99f[20]),
    .b(al_30e951fe[20]),
    .c(al_83614d40),
    .o({al_4182734,al_755dcbd4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c933ef2 (
    .a(al_e240f99f[21]),
    .b(al_30e951fe[21]),
    .c(al_4182734),
    .o({al_c006efbd,al_755dcbd4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_61814fa9 (
    .a(al_e240f99f[22]),
    .b(al_30e951fe[22]),
    .c(al_c006efbd),
    .o({al_49456793,al_755dcbd4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_94021f7e (
    .a(al_e240f99f[23]),
    .b(al_30e951fe[23]),
    .c(al_49456793),
    .o({al_e7a93f78,al_755dcbd4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9fe1b5e8 (
    .a(al_e240f99f[24]),
    .b(al_30e951fe[24]),
    .c(al_e7a93f78),
    .o({al_dd519345,al_755dcbd4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_339917e7 (
    .a(al_e240f99f[25]),
    .b(al_30e951fe[25]),
    .c(al_dd519345),
    .o({al_842cba6d,al_755dcbd4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_168be556 (
    .a(al_e240f99f[26]),
    .b(al_30e951fe[26]),
    .c(al_842cba6d),
    .o({al_bf0c2f5d,al_755dcbd4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de4c3c4 (
    .a(al_e240f99f[27]),
    .b(al_30e951fe[27]),
    .c(al_bf0c2f5d),
    .o({al_5059c5b1,al_755dcbd4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_622e61b3 (
    .a(al_e240f99f[28]),
    .b(al_30e951fe[28]),
    .c(al_5059c5b1),
    .o({al_cf4d3fd,al_755dcbd4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b49ecb6 (
    .a(al_e240f99f[29]),
    .b(al_30e951fe[29]),
    .c(al_cf4d3fd),
    .o({al_1df89094,al_755dcbd4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55beeada (
    .a(al_e240f99f[30]),
    .b(al_30e951fe[30]),
    .c(al_1df89094),
    .o({al_fdd90390,al_755dcbd4[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d3f533d6 (
    .a(al_e240f99f[31]),
    .b(al_30e951fe[31]),
    .c(al_fdd90390),
    .o({al_6e7e6fcf,al_755dcbd4[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_30bef3ee (
    .c(al_6e7e6fcf),
    .o({open_n59,al_755dcbd4[20]}));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_baf17d6e (
    .a(al_e8916352),
    .b(al_e240f99f[12]),
    .c(al_755dcbd4[0]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[12]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_7f15cc26 (
    .a(al_e8916352),
    .b(al_e240f99f[13]),
    .c(al_755dcbd4[1]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[13]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_d8d1a0a7 (
    .a(al_e8916352),
    .b(al_e240f99f[14]),
    .c(al_755dcbd4[2]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[14]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_651518d6 (
    .a(al_e8916352),
    .b(al_e240f99f[15]),
    .c(al_755dcbd4[3]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[15]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_9dea77b4 (
    .a(al_e8916352),
    .b(al_e240f99f[16]),
    .c(al_755dcbd4[4]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[16]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_b7a45d4b (
    .a(al_e8916352),
    .b(al_e240f99f[17]),
    .c(al_755dcbd4[5]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[17]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_605f5301 (
    .a(al_30e951fe[32]),
    .b(al_30e951fe[33]),
    .c(al_30e951fe[34]),
    .d(al_30e951fe[35]),
    .e(al_30e951fe[36]),
    .f(al_30e951fe[37]),
    .o(al_2daedad1));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_c2a59395 (
    .a(al_30e951fe[40]),
    .b(al_30e951fe[41]),
    .c(al_30e951fe[42]),
    .d(al_30e951fe[43]),
    .o(al_3b13cff4));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_301efbb2 (
    .a(al_2daedad1),
    .b(al_3b13cff4),
    .c(al_30e951fe[38]),
    .d(al_30e951fe[39]),
    .o(al_e8916352));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_cb4b63c8 (
    .a(al_e8916352),
    .b(al_e240f99f[18]),
    .c(al_755dcbd4[6]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[18]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_544bbf1 (
    .a(al_e8916352),
    .b(al_e240f99f[19]),
    .c(al_755dcbd4[7]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[19]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_929f6104 (
    .a(al_e8916352),
    .b(al_e240f99f[20]),
    .c(al_755dcbd4[8]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[20]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_9270245c (
    .a(al_e8916352),
    .b(al_e240f99f[21]),
    .c(al_755dcbd4[9]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[21]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_18b2a398 (
    .a(al_e8916352),
    .b(al_e240f99f[22]),
    .c(al_755dcbd4[10]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[22]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_1c9304e4 (
    .a(al_e8916352),
    .b(al_e240f99f[23]),
    .c(al_755dcbd4[11]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[23]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_749e687 (
    .a(al_e8916352),
    .b(al_e240f99f[24]),
    .c(al_755dcbd4[12]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[24]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_ca2b69b (
    .a(al_e8916352),
    .b(al_e240f99f[25]),
    .c(al_755dcbd4[13]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[25]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_62bbe168 (
    .a(al_e8916352),
    .b(al_e240f99f[26]),
    .c(al_755dcbd4[14]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[26]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_227ac8dd (
    .a(al_e8916352),
    .b(al_e240f99f[27]),
    .c(al_755dcbd4[15]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[27]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_862f1392 (
    .a(al_e8916352),
    .b(al_e240f99f[28]),
    .c(al_755dcbd4[16]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[28]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_165c84e4 (
    .a(al_e8916352),
    .b(al_e240f99f[29]),
    .c(al_755dcbd4[17]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[29]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_dc5f0eed (
    .a(al_e8916352),
    .b(al_e240f99f[30]),
    .c(al_755dcbd4[18]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[30]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcce4))
    al_f068bf18 (
    .a(al_e8916352),
    .b(al_e240f99f[31]),
    .c(al_755dcbd4[19]),
    .d(al_755dcbd4[20]),
    .o(al_abd7cd63[31]));
  AL_DFF_X al_9d5df6fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b0a2efb7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1c8da1e8[0]));
  AL_DFF_X al_4071744e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[11]));
  AL_DFF_X al_b40da1c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[12]));
  AL_DFF_X al_6fbbc63b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[13]));
  AL_DFF_X al_fec10209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[14]));
  AL_DFF_X al_4c5e75d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[15]));
  AL_DFF_X al_77c9ec96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[16]));
  AL_DFF_X al_2e4068f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[17]));
  AL_DFF_X al_81bace42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[18]));
  AL_DFF_X al_8714c1bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[19]));
  AL_DFF_X al_15285507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[20]));
  AL_DFF_X al_c960fc2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[21]));
  AL_DFF_X al_90bc04a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[22]));
  AL_DFF_X al_45f04ad5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[23]));
  AL_DFF_X al_ded55ebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[24]));
  AL_DFF_X al_26bdf5dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[25]));
  AL_DFF_X al_e06d55c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[26]));
  AL_DFF_X al_27df2608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[27]));
  AL_DFF_X al_2f1aec18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[28]));
  AL_DFF_X al_fd30384b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[29]));
  AL_DFF_X al_4c98587b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[30]));
  AL_DFF_X al_d5f3db29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[31]));
  AL_DFF_X al_3e359640 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[32]));
  AL_DFF_X al_b0423daa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[33]));
  AL_DFF_X al_74e767b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[34]));
  AL_DFF_X al_a195f5e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[35]));
  AL_DFF_X al_88fa2fd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[36]));
  AL_DFF_X al_1b90b50b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[37]));
  AL_DFF_X al_ad861fc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[38]));
  AL_DFF_X al_4478b361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[39]));
  AL_DFF_X al_737f8968 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[40]));
  AL_DFF_X al_2cc95497 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[41]));
  AL_DFF_X al_3f5c4fc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[42]));
  AL_DFF_X al_f9c20fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[8]));
  AL_DFF_X al_d3c76940 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[9]));
  AL_DFF_X al_c84c11e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[10]));
  AL_DFF_X al_293b13df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[11]));
  AL_DFF_X al_89a0c4c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[12]));
  AL_DFF_X al_29439f8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[13]));
  AL_DFF_X al_6954720d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[14]));
  AL_DFF_X al_ad11931a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[15]));
  AL_DFF_X al_4fb6ad44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[16]));
  AL_DFF_X al_d09e090c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[17]));
  AL_DFF_X al_8bdf081c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[0]));
  AL_DFF_X al_2127e46e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[18]));
  AL_DFF_X al_581460b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[19]));
  AL_DFF_X al_e59eb36d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[20]));
  AL_DFF_X al_2fa5500a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[21]));
  AL_DFF_X al_d65bf27f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[22]));
  AL_DFF_X al_690b5cef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[23]));
  AL_DFF_X al_4bdd3da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[24]));
  AL_DFF_X al_7e0ac317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[25]));
  AL_DFF_X al_3456c0bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[26]));
  AL_DFF_X al_5cc15d49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[27]));
  AL_DFF_X al_dad53c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[1]));
  AL_DFF_X al_cee402e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[28]));
  AL_DFF_X al_fd398974 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[29]));
  AL_DFF_X al_eae076a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[30]));
  AL_DFF_X al_f1df3b34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[31]));
  AL_DFF_X al_abf0ac53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[2]));
  AL_DFF_X al_66b0c258 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[3]));
  AL_DFF_X al_6c398f32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[4]));
  AL_DFF_X al_c034ca22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[5]));
  AL_DFF_X al_769956e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[6]));
  AL_DFF_X al_258252dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[7]));
  AL_DFF_X al_bf5c38f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[8]));
  AL_DFF_X al_74236897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[9]));
  AL_DFF_X al_be85bfc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[10]));
  AL_DFF_X al_8f8038fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[11]));
  AL_DFF_X al_f1bc7e23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[12]));
  AL_DFF_X al_726d2507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[13]));
  AL_DFF_X al_5a8cd6b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[14]));
  AL_DFF_X al_e39bc18a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[15]));
  AL_DFF_X al_a4f864a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[16]));
  AL_DFF_X al_e66b01d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[17]));
  AL_DFF_X al_50807c59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cc19a77c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[0]));
  AL_DFF_X al_a8640eee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[18]));
  AL_DFF_X al_479a297c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[19]));
  AL_DFF_X al_ed2f42cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[1]));
  AL_DFF_X al_c77bab5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[2]));
  AL_DFF_X al_e968a732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[3]));
  AL_DFF_X al_b6ba3a4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[4]));
  AL_DFF_X al_2fce49ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[5]));
  AL_DFF_X al_ec5c88b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[6]));
  AL_DFF_X al_f8d145a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    .INIT(16'hf731))
    al_d71568d (
    .a(al_3bd314e4[30]),
    .b(al_3bd314e4[31]),
    .c(al_83a08f3f[30]),
    .d(al_83a08f3f[31]),
    .o(al_e856fef8));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_4c9ec4fb (
    .a(al_2af03fa4),
    .b(al_b2d82920),
    .c(al_62013390),
    .d(al_e856fef8),
    .e(al_885349b2),
    .o(al_ebf67b92));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_cfdcda13 (
    .a(al_3bd314e4[38]),
    .b(al_3bd314e4[41]),
    .c(al_3bd314e4[43]),
    .d(al_3bd314e4[44]),
    .e(al_3bd314e4[46]),
    .f(al_3bd314e4[49]),
    .o(al_2ca9607b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_2add9bc5 (
    .a(al_3bd314e4[39]),
    .b(al_3bd314e4[40]),
    .c(al_3bd314e4[42]),
    .d(al_3bd314e4[45]),
    .o(al_13bec3a1));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_81b446c7 (
    .a(al_13bec3a1),
    .b(al_3bd314e4[32]),
    .c(al_3bd314e4[33]),
    .d(al_3bd314e4[34]),
    .e(al_3bd314e4[37]),
    .o(al_62013390));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_4296843c (
    .a(al_3bd314e4[35]),
    .b(al_3bd314e4[36]),
    .o(al_885349b2));
  AL_MAP_LUT4 #(
    .EQN("(A*(~(B)*C*~(D)+~(B)*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT(16'ha220))
    al_88dfe9af (
    .a(al_3bd314e4[30]),
    .b(al_3bd314e4[31]),
    .c(al_83a08f3f[30]),
    .d(al_83a08f3f[31]),
    .o(al_905b8225));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_8dff820c (
    .a(al_2af03fa4),
    .b(al_b2d82920),
    .c(al_62013390),
    .d(al_905b8225),
    .e(al_885349b2),
    .f(al_83a08f3f[30]),
    .o(al_89f2771a[30]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_507ef224 (
    .a(al_3bd314e4[55]),
    .b(al_3bd314e4[56]),
    .c(al_3bd314e4[58]),
    .d(al_3bd314e4[61]),
    .o(al_90792e1b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_a16a9bb5 (
    .a(al_2ca9607b),
    .b(al_90792e1b),
    .c(al_3bd314e4[51]),
    .d(al_3bd314e4[52]),
    .o(al_2af03fa4));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_9af2dddd (
    .a(al_3bd314e4[54]),
    .b(al_3bd314e4[57]),
    .c(al_3bd314e4[59]),
    .d(al_3bd314e4[60]),
    .o(al_9b8ff49a));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_8981c8e2 (
    .a(al_9b8ff49a),
    .b(al_3bd314e4[47]),
    .c(al_3bd314e4[48]),
    .d(al_3bd314e4[50]),
    .e(al_3bd314e4[53]),
    .o(al_b2d82920));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*A))"),
    .INIT(8'hc6))
    al_7c503c69 (
    .a(al_3bd314e4[30]),
    .b(al_3bd314e4[31]),
    .c(al_83a08f3f[30]),
    .o(al_3317fa82));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E*D*C*B*A))"),
    .INIT(64'h7fffffff00000000))
    al_f300627a (
    .a(al_2af03fa4),
    .b(al_b2d82920),
    .c(al_62013390),
    .d(al_3317fa82),
    .e(al_885349b2),
    .f(al_83a08f3f[31]),
    .o(al_89f2771a[31]));
  AL_DFF_X al_f4823322 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3da4ff6f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67f5b0b3[0]));
  AL_DFF_X al_d0b5d0bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[29]));
  AL_DFF_X al_6501b13d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[30]));
  AL_DFF_X al_ef9825f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[31]));
  AL_DFF_X al_2b73f5c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[32]));
  AL_DFF_X al_8eb770db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[33]));
  AL_DFF_X al_7b6ffac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[34]));
  AL_DFF_X al_9d18d894 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[35]));
  AL_DFF_X al_4d6f45d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[36]));
  AL_DFF_X al_638ccd8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[37]));
  AL_DFF_X al_10f6be35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[38]));
  AL_DFF_X al_92e646ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[39]));
  AL_DFF_X al_6d07d7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[40]));
  AL_DFF_X al_5cf08fb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[41]));
  AL_DFF_X al_3b5ceb01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[42]));
  AL_DFF_X al_43cfe69e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[43]));
  AL_DFF_X al_55fa205d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[44]));
  AL_DFF_X al_a51e3f0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[45]));
  AL_DFF_X al_cc73037d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[46]));
  AL_DFF_X al_3252fb45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[47]));
  AL_DFF_X al_2b0e150f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[48]));
  AL_DFF_X al_e6e3db5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[49]));
  AL_DFF_X al_17a6be0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[50]));
  AL_DFF_X al_a43099a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[51]));
  AL_DFF_X al_57e67c3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[52]));
  AL_DFF_X al_f08f3566 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[53]));
  AL_DFF_X al_964a5ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[54]));
  AL_DFF_X al_b190ee88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[55]));
  AL_DFF_X al_af6ce708 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[56]));
  AL_DFF_X al_785320fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[57]));
  AL_DFF_X al_48ca9fae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[58]));
  AL_DFF_X al_9cf96732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[59]));
  AL_DFF_X al_e3b7ef46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[60]));
  AL_DFF_X al_b4d44bea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[8]));
  AL_DFF_X al_4a2165bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[9]));
  AL_DFF_X al_de2727fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[10]));
  AL_DFF_X al_f1f71705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[11]));
  AL_DFF_X al_b81d9e59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[12]));
  AL_DFF_X al_eff51df1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[13]));
  AL_DFF_X al_15caecc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[14]));
  AL_DFF_X al_37b77fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[15]));
  AL_DFF_X al_a45082a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[16]));
  AL_DFF_X al_83c4c433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[17]));
  AL_DFF_X al_6faf62eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[0]));
  AL_DFF_X al_fcff1ea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[18]));
  AL_DFF_X al_2df0caf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[19]));
  AL_DFF_X al_7c4db8d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[20]));
  AL_DFF_X al_aad547ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[21]));
  AL_DFF_X al_e9321099 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[22]));
  AL_DFF_X al_17babbc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[23]));
  AL_DFF_X al_88e71fa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[24]));
  AL_DFF_X al_8bd27a00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[25]));
  AL_DFF_X al_f5cd7a87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[26]));
  AL_DFF_X al_e077ca3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[27]));
  AL_DFF_X al_af3f0e21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[1]));
  AL_DFF_X al_93861bd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[28]));
  AL_DFF_X al_7d029611 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[29]));
  AL_DFF_X al_8cb562a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_89f2771a[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[30]));
  AL_DFF_X al_4ed7d62b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_89f2771a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[31]));
  AL_DFF_X al_c55bc695 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[2]));
  AL_DFF_X al_5a7963d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[3]));
  AL_DFF_X al_896269e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[4]));
  AL_DFF_X al_afa1fbb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[5]));
  AL_DFF_X al_433bcd3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[6]));
  AL_DFF_X al_944b5435 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[7]));
  AL_DFF_X al_290f4151 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebf67b92),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b54c1014[0]));
  AL_DFF_X al_9cb2d599 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_33c3313d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b54c1014[1]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d6edf0c5 (
    .a(1'b0),
    .o({al_3b01c73c,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_504b6bae (
    .a(al_80a0f09e[11]),
    .b(al_e803eabe[11]),
    .c(al_3b01c73c),
    .o({al_5f9be50,al_ceb4d3af[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2838a311 (
    .a(al_80a0f09e[12]),
    .b(al_e803eabe[12]),
    .c(al_5f9be50),
    .o({al_c495520b,al_ceb4d3af[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_309339a4 (
    .a(al_80a0f09e[13]),
    .b(al_e803eabe[13]),
    .c(al_c495520b),
    .o({al_31fa6069,al_ceb4d3af[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_29176f29 (
    .a(al_80a0f09e[14]),
    .b(al_e803eabe[14]),
    .c(al_31fa6069),
    .o({al_add99006,al_ceb4d3af[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9cc5d94f (
    .a(al_80a0f09e[15]),
    .b(al_e803eabe[15]),
    .c(al_add99006),
    .o({al_3c7582f0,al_ceb4d3af[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8579bb6e (
    .a(al_80a0f09e[16]),
    .b(al_e803eabe[16]),
    .c(al_3c7582f0),
    .o({al_ad366bd4,al_ceb4d3af[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b67323c (
    .a(al_80a0f09e[17]),
    .b(al_e803eabe[17]),
    .c(al_ad366bd4),
    .o({al_435dca9c,al_ceb4d3af[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b986040e (
    .a(al_80a0f09e[18]),
    .b(al_e803eabe[18]),
    .c(al_435dca9c),
    .o({al_5689e405,al_ceb4d3af[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d264cd2b (
    .a(al_80a0f09e[19]),
    .b(al_e803eabe[19]),
    .c(al_5689e405),
    .o({al_af9115e4,al_ceb4d3af[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59f073a (
    .a(al_80a0f09e[20]),
    .b(al_e803eabe[20]),
    .c(al_af9115e4),
    .o({al_60435cbc,al_ceb4d3af[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f152d55 (
    .a(al_80a0f09e[21]),
    .b(al_e803eabe[21]),
    .c(al_60435cbc),
    .o({al_e0c9a948,al_ceb4d3af[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5343a940 (
    .a(al_80a0f09e[22]),
    .b(al_e803eabe[22]),
    .c(al_e0c9a948),
    .o({al_402ba912,al_ceb4d3af[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_510da646 (
    .a(al_80a0f09e[23]),
    .b(al_e803eabe[23]),
    .c(al_402ba912),
    .o({al_8caee7aa,al_ceb4d3af[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_681bfb5e (
    .a(al_80a0f09e[24]),
    .b(al_e803eabe[24]),
    .c(al_8caee7aa),
    .o({al_b7e03ff,al_ceb4d3af[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef1252c1 (
    .a(al_80a0f09e[25]),
    .b(al_e803eabe[25]),
    .c(al_b7e03ff),
    .o({al_74039666,al_ceb4d3af[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9e7ed8bb (
    .a(al_80a0f09e[26]),
    .b(al_e803eabe[26]),
    .c(al_74039666),
    .o({al_9da6bf97,al_ceb4d3af[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f71fe7b2 (
    .a(al_80a0f09e[27]),
    .b(al_e803eabe[27]),
    .c(al_9da6bf97),
    .o({al_23c46bef,al_ceb4d3af[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c561625e (
    .a(al_80a0f09e[28]),
    .b(al_e803eabe[28]),
    .c(al_23c46bef),
    .o({al_8c81e3ca,al_ceb4d3af[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45cb76dc (
    .a(al_80a0f09e[29]),
    .b(al_e803eabe[29]),
    .c(al_8c81e3ca),
    .o({al_f64316,al_ceb4d3af[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a1cf84a (
    .a(al_80a0f09e[30]),
    .b(al_e803eabe[30]),
    .c(al_f64316),
    .o({al_be55634f,al_ceb4d3af[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b26ad864 (
    .a(al_80a0f09e[31]),
    .b(al_e803eabe[31]),
    .c(al_be55634f),
    .o({al_631a2483,al_ceb4d3af[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f8bbbcd (
    .c(al_631a2483),
    .o({open_n65,al_ceb4d3af[21]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_51ebe859 (
    .a(al_e67fe640),
    .b(al_80a0f09e[11]),
    .c(al_ceb4d3af[0]),
    .o(al_cdad9264[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1614cf6c (
    .a(al_e67fe640),
    .b(al_80a0f09e[12]),
    .c(al_ceb4d3af[1]),
    .o(al_cdad9264[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_71fee9d (
    .a(al_e67fe640),
    .b(al_80a0f09e[13]),
    .c(al_ceb4d3af[2]),
    .o(al_cdad9264[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a5156781 (
    .a(al_e67fe640),
    .b(al_80a0f09e[14]),
    .c(al_ceb4d3af[3]),
    .o(al_cdad9264[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1aaf9798 (
    .a(al_e67fe640),
    .b(al_80a0f09e[15]),
    .c(al_ceb4d3af[4]),
    .o(al_cdad9264[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bc4f0586 (
    .a(al_e67fe640),
    .b(al_80a0f09e[16]),
    .c(al_ceb4d3af[5]),
    .o(al_cdad9264[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_69de076f (
    .a(al_e67fe640),
    .b(al_80a0f09e[17]),
    .c(al_ceb4d3af[6]),
    .o(al_cdad9264[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c72bf308 (
    .a(al_e67fe640),
    .b(al_80a0f09e[18]),
    .c(al_ceb4d3af[7]),
    .o(al_cdad9264[18]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b5a7a3f1 (
    .a(al_e803eabe[32]),
    .b(al_e803eabe[33]),
    .c(al_e803eabe[34]),
    .d(al_e803eabe[35]),
    .e(al_e803eabe[36]),
    .f(al_e803eabe[37]),
    .o(al_f8dbc1a1));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6b3ef705 (
    .a(al_e803eabe[40]),
    .b(al_e803eabe[41]),
    .c(al_e803eabe[42]),
    .d(al_ceb4d3af[21]),
    .o(al_ba13973b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_9eee0dc9 (
    .a(al_f8dbc1a1),
    .b(al_ba13973b),
    .c(al_e803eabe[38]),
    .d(al_e803eabe[39]),
    .o(al_e67fe640));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2330a9d (
    .a(al_e67fe640),
    .b(al_80a0f09e[19]),
    .c(al_ceb4d3af[8]),
    .o(al_cdad9264[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_16e19409 (
    .a(al_e67fe640),
    .b(al_80a0f09e[20]),
    .c(al_ceb4d3af[9]),
    .o(al_cdad9264[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e1ad6ee9 (
    .a(al_e67fe640),
    .b(al_80a0f09e[21]),
    .c(al_ceb4d3af[10]),
    .o(al_cdad9264[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b754c296 (
    .a(al_e67fe640),
    .b(al_80a0f09e[22]),
    .c(al_ceb4d3af[11]),
    .o(al_cdad9264[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_22254297 (
    .a(al_e67fe640),
    .b(al_80a0f09e[23]),
    .c(al_ceb4d3af[12]),
    .o(al_cdad9264[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1733a22f (
    .a(al_e67fe640),
    .b(al_80a0f09e[24]),
    .c(al_ceb4d3af[13]),
    .o(al_cdad9264[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d08110ed (
    .a(al_e67fe640),
    .b(al_80a0f09e[25]),
    .c(al_ceb4d3af[14]),
    .o(al_cdad9264[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_928b42b6 (
    .a(al_e67fe640),
    .b(al_80a0f09e[26]),
    .c(al_ceb4d3af[15]),
    .o(al_cdad9264[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_462139c4 (
    .a(al_e67fe640),
    .b(al_80a0f09e[27]),
    .c(al_ceb4d3af[16]),
    .o(al_cdad9264[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9c0350ac (
    .a(al_e67fe640),
    .b(al_80a0f09e[28]),
    .c(al_ceb4d3af[17]),
    .o(al_cdad9264[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_add5fc3f (
    .a(al_e67fe640),
    .b(al_80a0f09e[29]),
    .c(al_ceb4d3af[18]),
    .o(al_cdad9264[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e94977e (
    .a(al_e67fe640),
    .b(al_80a0f09e[30]),
    .c(al_ceb4d3af[19]),
    .o(al_cdad9264[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_58f6f719 (
    .a(al_e67fe640),
    .b(al_80a0f09e[31]),
    .c(al_ceb4d3af[20]),
    .o(al_cdad9264[31]));
  AL_DFF_X al_1c094ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c8da1e8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_acb3303d[0]));
  AL_DFF_X al_aad69b55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[10]));
  AL_DFF_X al_d5fc695 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[11]));
  AL_DFF_X al_9c7fa6d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[12]));
  AL_DFF_X al_2a9f2334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[13]));
  AL_DFF_X al_6e9cb2f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[14]));
  AL_DFF_X al_75f84619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[15]));
  AL_DFF_X al_77e56b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[16]));
  AL_DFF_X al_9495f3c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[17]));
  AL_DFF_X al_4160b8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[18]));
  AL_DFF_X al_80374bab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[19]));
  AL_DFF_X al_d4240dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[20]));
  AL_DFF_X al_58fc7f6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[21]));
  AL_DFF_X al_bf6c3422 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[22]));
  AL_DFF_X al_29644803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[23]));
  AL_DFF_X al_538903f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[24]));
  AL_DFF_X al_cb84a1ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[25]));
  AL_DFF_X al_bf40d6e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[26]));
  AL_DFF_X al_e67252ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[27]));
  AL_DFF_X al_e5dbf51e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[28]));
  AL_DFF_X al_5a0ab6bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[29]));
  AL_DFF_X al_29d9dc3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[30]));
  AL_DFF_X al_8bdebd35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[31]));
  AL_DFF_X al_5dc868c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[32]));
  AL_DFF_X al_7d00d0d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[33]));
  AL_DFF_X al_78cf7d7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[34]));
  AL_DFF_X al_4d829e30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[35]));
  AL_DFF_X al_c0ba87de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[36]));
  AL_DFF_X al_d25ae61b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[37]));
  AL_DFF_X al_6812a6ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[38]));
  AL_DFF_X al_39d0464e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[39]));
  AL_DFF_X al_7443e96f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[40]));
  AL_DFF_X al_c1f7e03e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[41]));
  AL_DFF_X al_ad0af11c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[8]));
  AL_DFF_X al_1e360c7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[9]));
  AL_DFF_X al_66d73fa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[10]));
  AL_DFF_X al_a72f1960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[11]));
  AL_DFF_X al_f9313079 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[12]));
  AL_DFF_X al_22b557f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[13]));
  AL_DFF_X al_dabe811f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[14]));
  AL_DFF_X al_e7dc64c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[15]));
  AL_DFF_X al_deac4ace (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[16]));
  AL_DFF_X al_abd30a62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[17]));
  AL_DFF_X al_9cbd4bf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[0]));
  AL_DFF_X al_ba76b98b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[18]));
  AL_DFF_X al_32b8ee78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[19]));
  AL_DFF_X al_81ec713c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[20]));
  AL_DFF_X al_e3177ad0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[21]));
  AL_DFF_X al_576615c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[22]));
  AL_DFF_X al_4643f5e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[23]));
  AL_DFF_X al_5595c4af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[24]));
  AL_DFF_X al_6f45a71c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[25]));
  AL_DFF_X al_51a6f581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[26]));
  AL_DFF_X al_41b20b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[27]));
  AL_DFF_X al_1455c68a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[1]));
  AL_DFF_X al_8aea6c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[28]));
  AL_DFF_X al_1ec12c43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[29]));
  AL_DFF_X al_1b984893 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[30]));
  AL_DFF_X al_ee695fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[31]));
  AL_DFF_X al_8fec86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[2]));
  AL_DFF_X al_52233176 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[3]));
  AL_DFF_X al_3a980319 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[4]));
  AL_DFF_X al_3707664f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[5]));
  AL_DFF_X al_466871e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[6]));
  AL_DFF_X al_3867c81e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[7]));
  AL_DFF_X al_99582d76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[8]));
  AL_DFF_X al_30eb1941 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[9]));
  AL_DFF_X al_2dd5f8e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[10]));
  AL_DFF_X al_84ec62a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[11]));
  AL_DFF_X al_1601700d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[12]));
  AL_DFF_X al_d75adf25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[13]));
  AL_DFF_X al_7191014d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[14]));
  AL_DFF_X al_2328cae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[15]));
  AL_DFF_X al_e53f998e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[16]));
  AL_DFF_X al_70840760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[17]));
  AL_DFF_X al_8004178b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e67fe640),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[0]));
  AL_DFF_X al_37f2080f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[18]));
  AL_DFF_X al_3e1a1112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[19]));
  AL_DFF_X al_d560510a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[20]));
  AL_DFF_X al_b08e1037 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[1]));
  AL_DFF_X al_b38d2529 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[2]));
  AL_DFF_X al_e7b53e70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[3]));
  AL_DFF_X al_61e5ffab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[4]));
  AL_DFF_X al_e072cf6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[5]));
  AL_DFF_X al_4ae4c2d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[6]));
  AL_DFF_X al_97bc4683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_649eda8a (
    .a(1'b0),
    .o({al_7f8fdeae,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e3f0e8ac (
    .a(al_98494645[10]),
    .b(al_753f5f88[10]),
    .c(al_7f8fdeae),
    .o({al_9d447f48,al_c706fd91[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5e6dd0a (
    .a(al_98494645[11]),
    .b(al_753f5f88[11]),
    .c(al_9d447f48),
    .o({al_56164bd3,al_c706fd91[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2c86c60 (
    .a(al_98494645[12]),
    .b(al_753f5f88[12]),
    .c(al_56164bd3),
    .o({al_f9511aee,al_c706fd91[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cabb207f (
    .a(al_98494645[13]),
    .b(al_753f5f88[13]),
    .c(al_f9511aee),
    .o({al_6a25f3ea,al_c706fd91[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47056f67 (
    .a(al_98494645[14]),
    .b(al_753f5f88[14]),
    .c(al_6a25f3ea),
    .o({al_abf34df7,al_c706fd91[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f79b43d7 (
    .a(al_98494645[15]),
    .b(al_753f5f88[15]),
    .c(al_abf34df7),
    .o({al_a6796ab,al_c706fd91[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_226d8e25 (
    .a(al_98494645[16]),
    .b(al_753f5f88[16]),
    .c(al_a6796ab),
    .o({al_59ba0f55,al_c706fd91[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_762a8eb3 (
    .a(al_98494645[17]),
    .b(al_753f5f88[17]),
    .c(al_59ba0f55),
    .o({al_92ed39a9,al_c706fd91[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f05c5980 (
    .a(al_98494645[18]),
    .b(al_753f5f88[18]),
    .c(al_92ed39a9),
    .o({al_c6dcc95e,al_c706fd91[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_371039af (
    .a(al_98494645[19]),
    .b(al_753f5f88[19]),
    .c(al_c6dcc95e),
    .o({al_1f87453b,al_c706fd91[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5d5a4ca (
    .a(al_98494645[20]),
    .b(al_753f5f88[20]),
    .c(al_1f87453b),
    .o({al_4c52cca8,al_c706fd91[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d6a73da1 (
    .a(al_98494645[21]),
    .b(al_753f5f88[21]),
    .c(al_4c52cca8),
    .o({al_bf05760,al_c706fd91[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a1aba8c (
    .a(al_98494645[22]),
    .b(al_753f5f88[22]),
    .c(al_bf05760),
    .o({al_ceb7552e,al_c706fd91[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a90f8b6d (
    .a(al_98494645[23]),
    .b(al_753f5f88[23]),
    .c(al_ceb7552e),
    .o({al_56dc547b,al_c706fd91[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_992de6af (
    .a(al_98494645[24]),
    .b(al_753f5f88[24]),
    .c(al_56dc547b),
    .o({al_cd3ff18,al_c706fd91[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d21abed (
    .a(al_98494645[25]),
    .b(al_753f5f88[25]),
    .c(al_cd3ff18),
    .o({al_cee7ade2,al_c706fd91[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cb0d8d2b (
    .a(al_98494645[26]),
    .b(al_753f5f88[26]),
    .c(al_cee7ade2),
    .o({al_afdea3b6,al_c706fd91[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fb01ef87 (
    .a(al_98494645[27]),
    .b(al_753f5f88[27]),
    .c(al_afdea3b6),
    .o({al_ed22eb5b,al_c706fd91[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27041c93 (
    .a(al_98494645[28]),
    .b(al_753f5f88[28]),
    .c(al_ed22eb5b),
    .o({al_7894a2ed,al_c706fd91[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2744a133 (
    .a(al_98494645[29]),
    .b(al_753f5f88[29]),
    .c(al_7894a2ed),
    .o({al_c319c1b9,al_c706fd91[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2449778a (
    .a(al_98494645[30]),
    .b(al_753f5f88[30]),
    .c(al_c319c1b9),
    .o({al_3111d364,al_c706fd91[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_262cbeb3 (
    .a(al_98494645[31]),
    .b(al_753f5f88[31]),
    .c(al_3111d364),
    .o({al_4e50336d,al_c706fd91[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e1e7a0e2 (
    .c(al_4e50336d),
    .o({open_n71,al_c706fd91[22]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bfe066ee (
    .a(al_c83520d8),
    .b(al_98494645[10]),
    .c(al_c706fd91[0]),
    .o(al_f7ed724c[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1ca3805 (
    .a(al_c83520d8),
    .b(al_98494645[11]),
    .c(al_c706fd91[1]),
    .o(al_f7ed724c[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_78abb849 (
    .a(al_c83520d8),
    .b(al_98494645[12]),
    .c(al_c706fd91[2]),
    .o(al_f7ed724c[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ecbefa1c (
    .a(al_c83520d8),
    .b(al_98494645[13]),
    .c(al_c706fd91[3]),
    .o(al_f7ed724c[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9150cabd (
    .a(al_c83520d8),
    .b(al_98494645[14]),
    .c(al_c706fd91[4]),
    .o(al_f7ed724c[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_281275b3 (
    .a(al_c83520d8),
    .b(al_98494645[15]),
    .c(al_c706fd91[5]),
    .o(al_f7ed724c[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_273bd6b0 (
    .a(al_c83520d8),
    .b(al_98494645[16]),
    .c(al_c706fd91[6]),
    .o(al_f7ed724c[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fc5850a5 (
    .a(al_c83520d8),
    .b(al_98494645[17]),
    .c(al_c706fd91[7]),
    .o(al_f7ed724c[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d5cbf9b2 (
    .a(al_c83520d8),
    .b(al_98494645[18]),
    .c(al_c706fd91[8]),
    .o(al_f7ed724c[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_18bb7064 (
    .a(al_c83520d8),
    .b(al_98494645[19]),
    .c(al_c706fd91[9]),
    .o(al_f7ed724c[19]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_26738965 (
    .a(al_753f5f88[36]),
    .b(al_753f5f88[37]),
    .c(al_753f5f88[38]),
    .d(al_753f5f88[39]),
    .e(al_753f5f88[40]),
    .f(al_753f5f88[41]),
    .o(al_99511a1d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_91b5a8e5 (
    .a(al_99511a1d),
    .b(al_753f5f88[32]),
    .c(al_753f5f88[33]),
    .d(al_753f5f88[34]),
    .e(al_753f5f88[35]),
    .f(al_c706fd91[22]),
    .o(al_c83520d8));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_71d60484 (
    .a(al_c83520d8),
    .b(al_98494645[20]),
    .c(al_c706fd91[10]),
    .o(al_f7ed724c[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6f4c0d76 (
    .a(al_c83520d8),
    .b(al_98494645[21]),
    .c(al_c706fd91[11]),
    .o(al_f7ed724c[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6dc50956 (
    .a(al_c83520d8),
    .b(al_98494645[22]),
    .c(al_c706fd91[12]),
    .o(al_f7ed724c[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9892f28c (
    .a(al_c83520d8),
    .b(al_98494645[23]),
    .c(al_c706fd91[13]),
    .o(al_f7ed724c[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3dd1295c (
    .a(al_c83520d8),
    .b(al_98494645[24]),
    .c(al_c706fd91[14]),
    .o(al_f7ed724c[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_15f56474 (
    .a(al_c83520d8),
    .b(al_98494645[25]),
    .c(al_c706fd91[15]),
    .o(al_f7ed724c[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_18f302d2 (
    .a(al_c83520d8),
    .b(al_98494645[26]),
    .c(al_c706fd91[16]),
    .o(al_f7ed724c[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c538154a (
    .a(al_c83520d8),
    .b(al_98494645[27]),
    .c(al_c706fd91[17]),
    .o(al_f7ed724c[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e08f281b (
    .a(al_c83520d8),
    .b(al_98494645[28]),
    .c(al_c706fd91[18]),
    .o(al_f7ed724c[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99561eae (
    .a(al_c83520d8),
    .b(al_98494645[29]),
    .c(al_c706fd91[19]),
    .o(al_f7ed724c[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_369dde19 (
    .a(al_c83520d8),
    .b(al_98494645[30]),
    .c(al_c706fd91[20]),
    .o(al_f7ed724c[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e402e97 (
    .a(al_c83520d8),
    .b(al_98494645[31]),
    .c(al_c706fd91[21]),
    .o(al_f7ed724c[31]));
  AL_DFF_X al_b8c97755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_acb3303d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14a1a59a[0]));
  AL_DFF_X al_1bad7c3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[9]));
  AL_DFF_X al_6f778f84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[10]));
  AL_DFF_X al_917e86c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[11]));
  AL_DFF_X al_aed909ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[12]));
  AL_DFF_X al_b4504b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[13]));
  AL_DFF_X al_fbf40054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[14]));
  AL_DFF_X al_6dfd5e83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[15]));
  AL_DFF_X al_350522b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[16]));
  AL_DFF_X al_b3143e5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[17]));
  AL_DFF_X al_bf2fa84f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[18]));
  AL_DFF_X al_bd4c7ccd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[19]));
  AL_DFF_X al_82438c15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[20]));
  AL_DFF_X al_3d4f4b3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[21]));
  AL_DFF_X al_e03d4811 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[22]));
  AL_DFF_X al_9a0fe6a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[23]));
  AL_DFF_X al_9feba60e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[24]));
  AL_DFF_X al_49108e80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[25]));
  AL_DFF_X al_8f1289f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[26]));
  AL_DFF_X al_57c4cf51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[27]));
  AL_DFF_X al_9c4d9923 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[28]));
  AL_DFF_X al_970d4407 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[29]));
  AL_DFF_X al_49b1e59f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[30]));
  AL_DFF_X al_ba224f5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[31]));
  AL_DFF_X al_caba6613 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[32]));
  AL_DFF_X al_e269d1b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[33]));
  AL_DFF_X al_be7dce89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[34]));
  AL_DFF_X al_ea140eef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[35]));
  AL_DFF_X al_4db0bbd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[36]));
  AL_DFF_X al_122e3941 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[37]));
  AL_DFF_X al_8611033a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[38]));
  AL_DFF_X al_dc02a858 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[39]));
  AL_DFF_X al_1ce9722b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[40]));
  AL_DFF_X al_9c2c2f1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[8]));
  AL_DFF_X al_c2f0ecf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[9]));
  AL_DFF_X al_13b58271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[10]));
  AL_DFF_X al_ab6c6990 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[11]));
  AL_DFF_X al_dbfc30f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[12]));
  AL_DFF_X al_c3f8f818 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[13]));
  AL_DFF_X al_e59ddad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[14]));
  AL_DFF_X al_5ea6ac44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[15]));
  AL_DFF_X al_5aac4542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[16]));
  AL_DFF_X al_e125a688 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[17]));
  AL_DFF_X al_e790fbae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[0]));
  AL_DFF_X al_b78716ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[18]));
  AL_DFF_X al_f2603864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[19]));
  AL_DFF_X al_58a3aee6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[20]));
  AL_DFF_X al_352316f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[21]));
  AL_DFF_X al_2434fe71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[22]));
  AL_DFF_X al_4a9b09dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[23]));
  AL_DFF_X al_a8a17df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[24]));
  AL_DFF_X al_b8293bc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[25]));
  AL_DFF_X al_8350ed20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[26]));
  AL_DFF_X al_bebe9a56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[27]));
  AL_DFF_X al_443d67af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[1]));
  AL_DFF_X al_aa0f98b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[28]));
  AL_DFF_X al_901194ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[29]));
  AL_DFF_X al_7f09e4bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[30]));
  AL_DFF_X al_560b977c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[31]));
  AL_DFF_X al_f9daadca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[2]));
  AL_DFF_X al_f017f428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[3]));
  AL_DFF_X al_ff5e7c13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[4]));
  AL_DFF_X al_88e32c30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[5]));
  AL_DFF_X al_11a98fcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[6]));
  AL_DFF_X al_55cc66bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[7]));
  AL_DFF_X al_ce3e18c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[8]));
  AL_DFF_X al_c9c77dec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[9]));
  AL_DFF_X al_5ac299e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[10]));
  AL_DFF_X al_80defe2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[11]));
  AL_DFF_X al_44cb480e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[12]));
  AL_DFF_X al_422ad121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[13]));
  AL_DFF_X al_bfd6e9bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[14]));
  AL_DFF_X al_9ef46c4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[15]));
  AL_DFF_X al_1305d5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[16]));
  AL_DFF_X al_5c640856 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[17]));
  AL_DFF_X al_fd0832b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c83520d8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[0]));
  AL_DFF_X al_b9bc2277 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[18]));
  AL_DFF_X al_2a7e92f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[19]));
  AL_DFF_X al_71832838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[20]));
  AL_DFF_X al_70a1cf96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[21]));
  AL_DFF_X al_4cfcba7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[1]));
  AL_DFF_X al_b817c0b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[2]));
  AL_DFF_X al_34478ebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[3]));
  AL_DFF_X al_3ced7650 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[4]));
  AL_DFF_X al_1ffcf69b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[5]));
  AL_DFF_X al_169b2f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[6]));
  AL_DFF_X al_33372a7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f00e13bb (
    .a(1'b0),
    .o({al_d6fc0fa3,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e8972cd (
    .a(al_bf34d64d[9]),
    .b(al_35594bd9[9]),
    .c(al_d6fc0fa3),
    .o({al_5b46bf26,al_abd8c6ec[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17f872e5 (
    .a(al_bf34d64d[10]),
    .b(al_35594bd9[10]),
    .c(al_5b46bf26),
    .o({al_5094d9fc,al_abd8c6ec[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d1dc7cb (
    .a(al_bf34d64d[11]),
    .b(al_35594bd9[11]),
    .c(al_5094d9fc),
    .o({al_94cd1325,al_abd8c6ec[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47bbfe54 (
    .a(al_bf34d64d[12]),
    .b(al_35594bd9[12]),
    .c(al_94cd1325),
    .o({al_b9861408,al_abd8c6ec[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2375fe1e (
    .a(al_bf34d64d[13]),
    .b(al_35594bd9[13]),
    .c(al_b9861408),
    .o({al_976c5f9d,al_abd8c6ec[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ad83c316 (
    .a(al_bf34d64d[14]),
    .b(al_35594bd9[14]),
    .c(al_976c5f9d),
    .o({al_e586ffc9,al_abd8c6ec[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33261058 (
    .a(al_bf34d64d[15]),
    .b(al_35594bd9[15]),
    .c(al_e586ffc9),
    .o({al_b45c14e1,al_abd8c6ec[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e017d9d (
    .a(al_bf34d64d[16]),
    .b(al_35594bd9[16]),
    .c(al_b45c14e1),
    .o({al_1b1dea64,al_abd8c6ec[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_326e0d2f (
    .a(al_bf34d64d[17]),
    .b(al_35594bd9[17]),
    .c(al_1b1dea64),
    .o({al_4188fe4e,al_abd8c6ec[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_370e757b (
    .a(al_bf34d64d[18]),
    .b(al_35594bd9[18]),
    .c(al_4188fe4e),
    .o({al_de74a82,al_abd8c6ec[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec70eca0 (
    .a(al_bf34d64d[19]),
    .b(al_35594bd9[19]),
    .c(al_de74a82),
    .o({al_632e424b,al_abd8c6ec[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2284d1fc (
    .a(al_bf34d64d[20]),
    .b(al_35594bd9[20]),
    .c(al_632e424b),
    .o({al_7fd8d148,al_abd8c6ec[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acce1c0 (
    .a(al_bf34d64d[21]),
    .b(al_35594bd9[21]),
    .c(al_7fd8d148),
    .o({al_6d674526,al_abd8c6ec[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a18ad069 (
    .a(al_bf34d64d[22]),
    .b(al_35594bd9[22]),
    .c(al_6d674526),
    .o({al_fdad78c8,al_abd8c6ec[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ecac0b66 (
    .a(al_bf34d64d[23]),
    .b(al_35594bd9[23]),
    .c(al_fdad78c8),
    .o({al_6620847d,al_abd8c6ec[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c654c13c (
    .a(al_bf34d64d[24]),
    .b(al_35594bd9[24]),
    .c(al_6620847d),
    .o({al_f4867e16,al_abd8c6ec[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7788f79c (
    .a(al_bf34d64d[25]),
    .b(al_35594bd9[25]),
    .c(al_f4867e16),
    .o({al_1bdf229b,al_abd8c6ec[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8424c54 (
    .a(al_bf34d64d[26]),
    .b(al_35594bd9[26]),
    .c(al_1bdf229b),
    .o({al_3e7ed8c8,al_abd8c6ec[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2b268755 (
    .a(al_bf34d64d[27]),
    .b(al_35594bd9[27]),
    .c(al_3e7ed8c8),
    .o({al_354fda56,al_abd8c6ec[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4a6524b8 (
    .a(al_bf34d64d[28]),
    .b(al_35594bd9[28]),
    .c(al_354fda56),
    .o({al_2f8d1c1e,al_abd8c6ec[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8bcea917 (
    .a(al_bf34d64d[29]),
    .b(al_35594bd9[29]),
    .c(al_2f8d1c1e),
    .o({al_57929d06,al_abd8c6ec[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37163518 (
    .a(al_bf34d64d[30]),
    .b(al_35594bd9[30]),
    .c(al_57929d06),
    .o({al_325baf0c,al_abd8c6ec[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fff85c4 (
    .a(al_bf34d64d[31]),
    .b(al_35594bd9[31]),
    .c(al_325baf0c),
    .o({al_9079498a,al_abd8c6ec[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_51708c60 (
    .c(al_9079498a),
    .o({open_n77,al_abd8c6ec[23]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f29beeba (
    .a(al_7715910d),
    .b(al_bf34d64d[10]),
    .c(al_abd8c6ec[1]),
    .o(al_96533024[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6a118cf0 (
    .a(al_7715910d),
    .b(al_bf34d64d[11]),
    .c(al_abd8c6ec[2]),
    .o(al_96533024[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cf292310 (
    .a(al_7715910d),
    .b(al_bf34d64d[12]),
    .c(al_abd8c6ec[3]),
    .o(al_96533024[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfde4b6b (
    .a(al_7715910d),
    .b(al_bf34d64d[13]),
    .c(al_abd8c6ec[4]),
    .o(al_96533024[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_10804e97 (
    .a(al_7715910d),
    .b(al_bf34d64d[14]),
    .c(al_abd8c6ec[5]),
    .o(al_96533024[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a9786286 (
    .a(al_7715910d),
    .b(al_bf34d64d[15]),
    .c(al_abd8c6ec[6]),
    .o(al_96533024[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_52b72919 (
    .a(al_7715910d),
    .b(al_bf34d64d[16]),
    .c(al_abd8c6ec[7]),
    .o(al_96533024[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dabf5e16 (
    .a(al_7715910d),
    .b(al_bf34d64d[17]),
    .c(al_abd8c6ec[8]),
    .o(al_96533024[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da5d7bdf (
    .a(al_7715910d),
    .b(al_bf34d64d[18]),
    .c(al_abd8c6ec[9]),
    .o(al_96533024[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a28ee61b (
    .a(al_7715910d),
    .b(al_bf34d64d[19]),
    .c(al_abd8c6ec[10]),
    .o(al_96533024[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_146b2ad7 (
    .a(al_7715910d),
    .b(al_bf34d64d[20]),
    .c(al_abd8c6ec[11]),
    .o(al_96533024[20]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6cf4fc6c (
    .a(al_35594bd9[36]),
    .b(al_35594bd9[37]),
    .c(al_35594bd9[38]),
    .d(al_35594bd9[39]),
    .e(al_35594bd9[40]),
    .f(al_abd8c6ec[23]),
    .o(al_d2dbac27));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_6d1e3807 (
    .a(al_d2dbac27),
    .b(al_35594bd9[32]),
    .c(al_35594bd9[33]),
    .d(al_35594bd9[34]),
    .e(al_35594bd9[35]),
    .o(al_7715910d));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_43183a47 (
    .a(al_7715910d),
    .b(al_bf34d64d[21]),
    .c(al_abd8c6ec[12]),
    .o(al_96533024[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_67ad3d73 (
    .a(al_7715910d),
    .b(al_bf34d64d[22]),
    .c(al_abd8c6ec[13]),
    .o(al_96533024[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_43c3758d (
    .a(al_7715910d),
    .b(al_bf34d64d[23]),
    .c(al_abd8c6ec[14]),
    .o(al_96533024[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9619ffa (
    .a(al_7715910d),
    .b(al_bf34d64d[24]),
    .c(al_abd8c6ec[15]),
    .o(al_96533024[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c8755677 (
    .a(al_7715910d),
    .b(al_bf34d64d[25]),
    .c(al_abd8c6ec[16]),
    .o(al_96533024[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_15a71cc6 (
    .a(al_7715910d),
    .b(al_bf34d64d[26]),
    .c(al_abd8c6ec[17]),
    .o(al_96533024[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_85d5f343 (
    .a(al_7715910d),
    .b(al_bf34d64d[27]),
    .c(al_abd8c6ec[18]),
    .o(al_96533024[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfe9fd59 (
    .a(al_7715910d),
    .b(al_bf34d64d[28]),
    .c(al_abd8c6ec[19]),
    .o(al_96533024[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f01e5bc (
    .a(al_7715910d),
    .b(al_bf34d64d[29]),
    .c(al_abd8c6ec[20]),
    .o(al_96533024[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4c47521 (
    .a(al_7715910d),
    .b(al_bf34d64d[30]),
    .c(al_abd8c6ec[21]),
    .o(al_96533024[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b1a091eb (
    .a(al_7715910d),
    .b(al_bf34d64d[31]),
    .c(al_abd8c6ec[22]),
    .o(al_96533024[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b8a3d57f (
    .a(al_7715910d),
    .b(al_bf34d64d[9]),
    .c(al_abd8c6ec[0]),
    .o(al_96533024[9]));
  AL_DFF_X al_f66e1479 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14a1a59a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_21143207[0]));
  AL_DFF_X al_3e3b493b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[8]));
  AL_DFF_X al_1bd47a66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[9]));
  AL_DFF_X al_93223d64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[10]));
  AL_DFF_X al_b1e7de9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[11]));
  AL_DFF_X al_878fa54b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[12]));
  AL_DFF_X al_906c63e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[13]));
  AL_DFF_X al_ec61ff37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[14]));
  AL_DFF_X al_4c3558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[15]));
  AL_DFF_X al_89fadf24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[16]));
  AL_DFF_X al_b5d783a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[17]));
  AL_DFF_X al_ba4c82e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[18]));
  AL_DFF_X al_636eb843 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[19]));
  AL_DFF_X al_5672314d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[20]));
  AL_DFF_X al_3708b4aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[21]));
  AL_DFF_X al_1a14e6f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[22]));
  AL_DFF_X al_2953eb04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[23]));
  AL_DFF_X al_a31aaaf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[24]));
  AL_DFF_X al_bede1366 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[25]));
  AL_DFF_X al_b2e1fd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[26]));
  AL_DFF_X al_5946d8fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[27]));
  AL_DFF_X al_669887e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[28]));
  AL_DFF_X al_eed4127c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[29]));
  AL_DFF_X al_2906c568 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[30]));
  AL_DFF_X al_3ab403da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[31]));
  AL_DFF_X al_b7cedbe3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[32]));
  AL_DFF_X al_a8a427b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[33]));
  AL_DFF_X al_bc10962b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[34]));
  AL_DFF_X al_51c8b1cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[35]));
  AL_DFF_X al_3c1bd03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[36]));
  AL_DFF_X al_97c3ce00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[37]));
  AL_DFF_X al_f88eb3ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[38]));
  AL_DFF_X al_5aaedb4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[39]));
  AL_DFF_X al_9a7849ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[8]));
  AL_DFF_X al_6eeb394a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[9]));
  AL_DFF_X al_642c2710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[10]));
  AL_DFF_X al_f5734ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[11]));
  AL_DFF_X al_2fd7def (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[12]));
  AL_DFF_X al_61826c3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[13]));
  AL_DFF_X al_ebc885e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[14]));
  AL_DFF_X al_654d7630 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[15]));
  AL_DFF_X al_42ba68ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[16]));
  AL_DFF_X al_cb8e6d7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[17]));
  AL_DFF_X al_904222ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[0]));
  AL_DFF_X al_902523b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[18]));
  AL_DFF_X al_a152f96b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[19]));
  AL_DFF_X al_e783dbc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[20]));
  AL_DFF_X al_12c4b239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[21]));
  AL_DFF_X al_c986b495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[22]));
  AL_DFF_X al_a7b8dfbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[23]));
  AL_DFF_X al_7a2781e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[24]));
  AL_DFF_X al_aae3d656 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[25]));
  AL_DFF_X al_3e3a5494 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[26]));
  AL_DFF_X al_6ea11ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[27]));
  AL_DFF_X al_1a4cb7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[1]));
  AL_DFF_X al_cf76b977 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[28]));
  AL_DFF_X al_96df0728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[29]));
  AL_DFF_X al_688a3213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[30]));
  AL_DFF_X al_474f4d26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[31]));
  AL_DFF_X al_c5c3843f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[2]));
  AL_DFF_X al_dd27dfcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[3]));
  AL_DFF_X al_f4ddc2f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[4]));
  AL_DFF_X al_1bb5d678 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[5]));
  AL_DFF_X al_c3e4d2d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[6]));
  AL_DFF_X al_aec44769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[7]));
  AL_DFF_X al_d7924fdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[8]));
  AL_DFF_X al_13943ca8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[9]));
  AL_DFF_X al_3121d73f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[10]));
  AL_DFF_X al_8f17eb61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[11]));
  AL_DFF_X al_a1ef3bd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[12]));
  AL_DFF_X al_af8a903b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[13]));
  AL_DFF_X al_772b7806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[14]));
  AL_DFF_X al_cd8f8f12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[15]));
  AL_DFF_X al_6cbe6158 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[16]));
  AL_DFF_X al_c7b21531 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[17]));
  AL_DFF_X al_460715fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7715910d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[0]));
  AL_DFF_X al_38d6e179 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[18]));
  AL_DFF_X al_60fe0a64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[19]));
  AL_DFF_X al_eaa5b1be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[20]));
  AL_DFF_X al_6609171e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[21]));
  AL_DFF_X al_76c593f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[22]));
  AL_DFF_X al_36a85cdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[1]));
  AL_DFF_X al_775775aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[2]));
  AL_DFF_X al_f0fae96b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[3]));
  AL_DFF_X al_851177b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[4]));
  AL_DFF_X al_7bf7fe43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[5]));
  AL_DFF_X al_5c587394 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[6]));
  AL_DFF_X al_22a47df5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ae71dfc7 (
    .a(1'b0),
    .o({al_f486a09d,open_n80}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b49808c (
    .a(al_f0f43754[8]),
    .b(al_f2bb4ec4[8]),
    .c(al_f486a09d),
    .o({al_bee033d9,al_801f6a4a[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d96fba64 (
    .a(al_f0f43754[9]),
    .b(al_f2bb4ec4[9]),
    .c(al_bee033d9),
    .o({al_a60df36b,al_801f6a4a[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eaf4f230 (
    .a(al_f0f43754[10]),
    .b(al_f2bb4ec4[10]),
    .c(al_a60df36b),
    .o({al_aa119f92,al_801f6a4a[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f66536f4 (
    .a(al_f0f43754[11]),
    .b(al_f2bb4ec4[11]),
    .c(al_aa119f92),
    .o({al_ced042bc,al_801f6a4a[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cd87d517 (
    .a(al_f0f43754[12]),
    .b(al_f2bb4ec4[12]),
    .c(al_ced042bc),
    .o({al_9de12621,al_801f6a4a[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a462211 (
    .a(al_f0f43754[13]),
    .b(al_f2bb4ec4[13]),
    .c(al_9de12621),
    .o({al_c6d35f30,al_801f6a4a[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_64593f54 (
    .a(al_f0f43754[14]),
    .b(al_f2bb4ec4[14]),
    .c(al_c6d35f30),
    .o({al_41de2ced,al_801f6a4a[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f875cb (
    .a(al_f0f43754[15]),
    .b(al_f2bb4ec4[15]),
    .c(al_41de2ced),
    .o({al_a4baa375,al_801f6a4a[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc86ab10 (
    .a(al_f0f43754[16]),
    .b(al_f2bb4ec4[16]),
    .c(al_a4baa375),
    .o({al_7d7301fd,al_801f6a4a[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e71fd686 (
    .a(al_f0f43754[17]),
    .b(al_f2bb4ec4[17]),
    .c(al_7d7301fd),
    .o({al_f804f442,al_801f6a4a[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d119fc0d (
    .a(al_f0f43754[18]),
    .b(al_f2bb4ec4[18]),
    .c(al_f804f442),
    .o({al_fa20e924,al_801f6a4a[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_df81cd21 (
    .a(al_f0f43754[19]),
    .b(al_f2bb4ec4[19]),
    .c(al_fa20e924),
    .o({al_75df31c,al_801f6a4a[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72a296c2 (
    .a(al_f0f43754[20]),
    .b(al_f2bb4ec4[20]),
    .c(al_75df31c),
    .o({al_fb6c6a88,al_801f6a4a[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_502880a5 (
    .a(al_f0f43754[21]),
    .b(al_f2bb4ec4[21]),
    .c(al_fb6c6a88),
    .o({al_6a47eaf1,al_801f6a4a[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d3245e45 (
    .a(al_f0f43754[22]),
    .b(al_f2bb4ec4[22]),
    .c(al_6a47eaf1),
    .o({al_ef2cb93b,al_801f6a4a[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e616607 (
    .a(al_f0f43754[23]),
    .b(al_f2bb4ec4[23]),
    .c(al_ef2cb93b),
    .o({al_7c6e81bc,al_801f6a4a[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9e0ee99 (
    .a(al_f0f43754[24]),
    .b(al_f2bb4ec4[24]),
    .c(al_7c6e81bc),
    .o({al_820ba18b,al_801f6a4a[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_75569f3c (
    .a(al_f0f43754[25]),
    .b(al_f2bb4ec4[25]),
    .c(al_820ba18b),
    .o({al_90eca21f,al_801f6a4a[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7520c3fb (
    .a(al_f0f43754[26]),
    .b(al_f2bb4ec4[26]),
    .c(al_90eca21f),
    .o({al_14135fe,al_801f6a4a[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8df74e6c (
    .a(al_f0f43754[27]),
    .b(al_f2bb4ec4[27]),
    .c(al_14135fe),
    .o({al_278fc7b9,al_801f6a4a[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed06cb72 (
    .a(al_f0f43754[28]),
    .b(al_f2bb4ec4[28]),
    .c(al_278fc7b9),
    .o({al_78f968d6,al_801f6a4a[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_208e0aef (
    .a(al_f0f43754[29]),
    .b(al_f2bb4ec4[29]),
    .c(al_78f968d6),
    .o({al_6cb6cc70,al_801f6a4a[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_63ab56df (
    .a(al_f0f43754[30]),
    .b(al_f2bb4ec4[30]),
    .c(al_6cb6cc70),
    .o({al_5bfcf8ca,al_801f6a4a[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c90ccf3 (
    .a(al_f0f43754[31]),
    .b(al_f2bb4ec4[31]),
    .c(al_5bfcf8ca),
    .o({al_7777e58e,al_801f6a4a[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_528a8d0c (
    .c(al_7777e58e),
    .o({open_n83,al_801f6a4a[24]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ec0d9fc2 (
    .a(al_665b7858),
    .b(al_f0f43754[10]),
    .c(al_801f6a4a[2]),
    .o(al_e60d8647[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c89256c (
    .a(al_665b7858),
    .b(al_f0f43754[11]),
    .c(al_801f6a4a[3]),
    .o(al_e60d8647[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_20d40a82 (
    .a(al_665b7858),
    .b(al_f0f43754[12]),
    .c(al_801f6a4a[4]),
    .o(al_e60d8647[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d8154562 (
    .a(al_665b7858),
    .b(al_f0f43754[13]),
    .c(al_801f6a4a[5]),
    .o(al_e60d8647[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_94a67f78 (
    .a(al_665b7858),
    .b(al_f0f43754[14]),
    .c(al_801f6a4a[6]),
    .o(al_e60d8647[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8ec18da0 (
    .a(al_665b7858),
    .b(al_f0f43754[15]),
    .c(al_801f6a4a[7]),
    .o(al_e60d8647[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6ae98376 (
    .a(al_665b7858),
    .b(al_f0f43754[16]),
    .c(al_801f6a4a[8]),
    .o(al_e60d8647[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c41b103d (
    .a(al_665b7858),
    .b(al_f0f43754[17]),
    .c(al_801f6a4a[9]),
    .o(al_e60d8647[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f9441d24 (
    .a(al_665b7858),
    .b(al_f0f43754[18]),
    .c(al_801f6a4a[10]),
    .o(al_e60d8647[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e90b325a (
    .a(al_665b7858),
    .b(al_f0f43754[19]),
    .c(al_801f6a4a[11]),
    .o(al_e60d8647[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f477e3c5 (
    .a(al_665b7858),
    .b(al_f0f43754[20]),
    .c(al_801f6a4a[12]),
    .o(al_e60d8647[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b9554dc4 (
    .a(al_665b7858),
    .b(al_f0f43754[21]),
    .c(al_801f6a4a[13]),
    .o(al_e60d8647[21]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_bcf7dcb6 (
    .a(al_f2bb4ec4[34]),
    .b(al_f2bb4ec4[35]),
    .c(al_f2bb4ec4[36]),
    .d(al_f2bb4ec4[37]),
    .e(al_f2bb4ec4[38]),
    .f(al_f2bb4ec4[39]),
    .o(al_ce2d0e53));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_922c9aa2 (
    .a(al_ce2d0e53),
    .b(al_f2bb4ec4[32]),
    .c(al_f2bb4ec4[33]),
    .d(al_801f6a4a[24]),
    .o(al_665b7858));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_413db73c (
    .a(al_665b7858),
    .b(al_f0f43754[22]),
    .c(al_801f6a4a[14]),
    .o(al_e60d8647[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0a44916 (
    .a(al_665b7858),
    .b(al_f0f43754[23]),
    .c(al_801f6a4a[15]),
    .o(al_e60d8647[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2fbc7b03 (
    .a(al_665b7858),
    .b(al_f0f43754[24]),
    .c(al_801f6a4a[16]),
    .o(al_e60d8647[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d796eadb (
    .a(al_665b7858),
    .b(al_f0f43754[25]),
    .c(al_801f6a4a[17]),
    .o(al_e60d8647[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4f8857c (
    .a(al_665b7858),
    .b(al_f0f43754[26]),
    .c(al_801f6a4a[18]),
    .o(al_e60d8647[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e6253bca (
    .a(al_665b7858),
    .b(al_f0f43754[27]),
    .c(al_801f6a4a[19]),
    .o(al_e60d8647[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c9732bef (
    .a(al_665b7858),
    .b(al_f0f43754[28]),
    .c(al_801f6a4a[20]),
    .o(al_e60d8647[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1491d4b7 (
    .a(al_665b7858),
    .b(al_f0f43754[29]),
    .c(al_801f6a4a[21]),
    .o(al_e60d8647[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9c82427f (
    .a(al_665b7858),
    .b(al_f0f43754[30]),
    .c(al_801f6a4a[22]),
    .o(al_e60d8647[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_47cb7671 (
    .a(al_665b7858),
    .b(al_f0f43754[31]),
    .c(al_801f6a4a[23]),
    .o(al_e60d8647[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_131b00fa (
    .a(al_665b7858),
    .b(al_f0f43754[8]),
    .c(al_801f6a4a[0]),
    .o(al_e60d8647[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_675e87c2 (
    .a(al_665b7858),
    .b(al_f0f43754[9]),
    .c(al_801f6a4a[1]),
    .o(al_e60d8647[9]));
  AL_DFF_X al_87358168 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_21143207[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e0dc7e9e[0]));
  AL_DFF_X al_d29dd6bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[8]));
  AL_DFF_X al_a288c327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[9]));
  AL_DFF_X al_6c67fd46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[10]));
  AL_DFF_X al_d8e0999a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[11]));
  AL_DFF_X al_62b4b794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[12]));
  AL_DFF_X al_1ac6a7f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[13]));
  AL_DFF_X al_b7561573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[14]));
  AL_DFF_X al_d117c4b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[15]));
  AL_DFF_X al_6ef3e2bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[16]));
  AL_DFF_X al_8a3809d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[17]));
  AL_DFF_X al_69711203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[18]));
  AL_DFF_X al_10aaaab0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[19]));
  AL_DFF_X al_4b859408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[20]));
  AL_DFF_X al_e14bc755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[21]));
  AL_DFF_X al_6527d3c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[22]));
  AL_DFF_X al_444b851f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[23]));
  AL_DFF_X al_e312d94f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[24]));
  AL_DFF_X al_f539dba2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[25]));
  AL_DFF_X al_f50f81ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[26]));
  AL_DFF_X al_59ecc5d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[27]));
  AL_DFF_X al_c3a6f296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[28]));
  AL_DFF_X al_fd8973ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[29]));
  AL_DFF_X al_ce9d9527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[30]));
  AL_DFF_X al_169f74c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[31]));
  AL_DFF_X al_6af3b830 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[32]));
  AL_DFF_X al_e9563b2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[33]));
  AL_DFF_X al_b4aa1ef4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[34]));
  AL_DFF_X al_1eddd24d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[35]));
  AL_DFF_X al_4cfb845 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[36]));
  AL_DFF_X al_96cdb566 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[37]));
  AL_DFF_X al_6ef0a018 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[38]));
  AL_DFF_X al_78620cd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[7]));
  AL_DFF_X al_6f93fd80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[8]));
  AL_DFF_X al_c99b16e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[9]));
  AL_DFF_X al_d5c10c50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[10]));
  AL_DFF_X al_5e81c9a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[11]));
  AL_DFF_X al_bf1169fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[12]));
  AL_DFF_X al_28d8c1b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[13]));
  AL_DFF_X al_ec3e6e83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[14]));
  AL_DFF_X al_f2062cec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[15]));
  AL_DFF_X al_a3afe68d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[16]));
  AL_DFF_X al_ec380358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[17]));
  AL_DFF_X al_f8e94199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[0]));
  AL_DFF_X al_f3f9c4d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[18]));
  AL_DFF_X al_6c0d985e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[19]));
  AL_DFF_X al_dfd344ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[20]));
  AL_DFF_X al_3c3daa43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[21]));
  AL_DFF_X al_7ffafa27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[22]));
  AL_DFF_X al_8d7046e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[23]));
  AL_DFF_X al_3df49cc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[24]));
  AL_DFF_X al_78653f90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[25]));
  AL_DFF_X al_5b757883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[26]));
  AL_DFF_X al_cce245e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[27]));
  AL_DFF_X al_7d132e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[1]));
  AL_DFF_X al_34ce0bbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[28]));
  AL_DFF_X al_2677c5b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[29]));
  AL_DFF_X al_232ad16b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[30]));
  AL_DFF_X al_7f25f5cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[31]));
  AL_DFF_X al_affd94a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[2]));
  AL_DFF_X al_f7d9f7e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[3]));
  AL_DFF_X al_f942d56e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[4]));
  AL_DFF_X al_935b35d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[5]));
  AL_DFF_X al_a30094fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[6]));
  AL_DFF_X al_2f9d854b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[7]));
  AL_DFF_X al_cb6e6a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[8]));
  AL_DFF_X al_fb2ced0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[9]));
  AL_DFF_X al_2967b583 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[10]));
  AL_DFF_X al_de9dea44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[11]));
  AL_DFF_X al_cf23a99c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[12]));
  AL_DFF_X al_8493f479 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[13]));
  AL_DFF_X al_60181410 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[14]));
  AL_DFF_X al_80c061bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[15]));
  AL_DFF_X al_d1b0ef37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[16]));
  AL_DFF_X al_9ce13146 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[17]));
  AL_DFF_X al_94085238 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_665b7858),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[0]));
  AL_DFF_X al_696af070 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[18]));
  AL_DFF_X al_5c3ad2bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[19]));
  AL_DFF_X al_8018de15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[20]));
  AL_DFF_X al_1bcdffa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[21]));
  AL_DFF_X al_ed3d0137 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[22]));
  AL_DFF_X al_599f4a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[23]));
  AL_DFF_X al_29f6d41f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[1]));
  AL_DFF_X al_6aa8574b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[2]));
  AL_DFF_X al_d58fa4fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[3]));
  AL_DFF_X al_3019f739 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[4]));
  AL_DFF_X al_57be8bae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[5]));
  AL_DFF_X al_dbb0a998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[6]));
  AL_DFF_X al_44c8a552 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_8ec5f588 (
    .a(1'b0),
    .o({al_3d0d887e,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b150ed4 (
    .a(al_86280a69[7]),
    .b(al_3029c49a[7]),
    .c(al_3d0d887e),
    .o({al_f44c949b,al_591ecc80[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9dc9e38f (
    .a(al_86280a69[8]),
    .b(al_3029c49a[8]),
    .c(al_f44c949b),
    .o({al_394ce23b,al_591ecc80[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_69949589 (
    .a(al_86280a69[9]),
    .b(al_3029c49a[9]),
    .c(al_394ce23b),
    .o({al_354fae1f,al_591ecc80[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e08dff4f (
    .a(al_86280a69[10]),
    .b(al_3029c49a[10]),
    .c(al_354fae1f),
    .o({al_89af750e,al_591ecc80[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e3e1db98 (
    .a(al_86280a69[11]),
    .b(al_3029c49a[11]),
    .c(al_89af750e),
    .o({al_8cf6cbd4,al_591ecc80[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_383abf3e (
    .a(al_86280a69[12]),
    .b(al_3029c49a[12]),
    .c(al_8cf6cbd4),
    .o({al_32030ed2,al_591ecc80[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_561806c6 (
    .a(al_86280a69[13]),
    .b(al_3029c49a[13]),
    .c(al_32030ed2),
    .o({al_5875f740,al_591ecc80[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_82ecb0d8 (
    .a(al_86280a69[14]),
    .b(al_3029c49a[14]),
    .c(al_5875f740),
    .o({al_7cb5ff51,al_591ecc80[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_274cc367 (
    .a(al_86280a69[15]),
    .b(al_3029c49a[15]),
    .c(al_7cb5ff51),
    .o({al_ee0cbe48,al_591ecc80[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88c06b23 (
    .a(al_86280a69[16]),
    .b(al_3029c49a[16]),
    .c(al_ee0cbe48),
    .o({al_b4749ad8,al_591ecc80[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3784d2 (
    .a(al_86280a69[17]),
    .b(al_3029c49a[17]),
    .c(al_b4749ad8),
    .o({al_dc8ef999,al_591ecc80[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e344ff48 (
    .a(al_86280a69[18]),
    .b(al_3029c49a[18]),
    .c(al_dc8ef999),
    .o({al_500654bb,al_591ecc80[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_568b2ece (
    .a(al_86280a69[19]),
    .b(al_3029c49a[19]),
    .c(al_500654bb),
    .o({al_62272aaf,al_591ecc80[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce568604 (
    .a(al_86280a69[20]),
    .b(al_3029c49a[20]),
    .c(al_62272aaf),
    .o({al_2f455704,al_591ecc80[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d80782ec (
    .a(al_86280a69[21]),
    .b(al_3029c49a[21]),
    .c(al_2f455704),
    .o({al_b7b82cb6,al_591ecc80[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8eb3be72 (
    .a(al_86280a69[22]),
    .b(al_3029c49a[22]),
    .c(al_b7b82cb6),
    .o({al_7375cfb0,al_591ecc80[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b7ebbb (
    .a(al_86280a69[23]),
    .b(al_3029c49a[23]),
    .c(al_7375cfb0),
    .o({al_c78e76e7,al_591ecc80[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a2590dc7 (
    .a(al_86280a69[24]),
    .b(al_3029c49a[24]),
    .c(al_c78e76e7),
    .o({al_ef33e959,al_591ecc80[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33ab491 (
    .a(al_86280a69[25]),
    .b(al_3029c49a[25]),
    .c(al_ef33e959),
    .o({al_6387fe,al_591ecc80[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e1a45f73 (
    .a(al_86280a69[26]),
    .b(al_3029c49a[26]),
    .c(al_6387fe),
    .o({al_25d9aae7,al_591ecc80[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_44052f24 (
    .a(al_86280a69[27]),
    .b(al_3029c49a[27]),
    .c(al_25d9aae7),
    .o({al_9233bdf0,al_591ecc80[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_753c5315 (
    .a(al_86280a69[28]),
    .b(al_3029c49a[28]),
    .c(al_9233bdf0),
    .o({al_cee8b982,al_591ecc80[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f0c68d81 (
    .a(al_86280a69[29]),
    .b(al_3029c49a[29]),
    .c(al_cee8b982),
    .o({al_c5ec6219,al_591ecc80[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f989d1cc (
    .a(al_86280a69[30]),
    .b(al_3029c49a[30]),
    .c(al_c5ec6219),
    .o({al_ae24ecf8,al_591ecc80[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6973685b (
    .a(al_86280a69[31]),
    .b(al_3029c49a[31]),
    .c(al_ae24ecf8),
    .o({al_72ba4be2,al_591ecc80[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1cea3bfa (
    .c(al_72ba4be2),
    .o({open_n89,al_591ecc80[25]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_63cdce2d (
    .a(al_2878e2ee),
    .b(al_86280a69[10]),
    .c(al_591ecc80[3]),
    .o(al_f78b30ce[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a580bb7e (
    .a(al_2878e2ee),
    .b(al_86280a69[11]),
    .c(al_591ecc80[4]),
    .o(al_f78b30ce[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_61740b7b (
    .a(al_2878e2ee),
    .b(al_86280a69[12]),
    .c(al_591ecc80[5]),
    .o(al_f78b30ce[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d12ca8de (
    .a(al_2878e2ee),
    .b(al_86280a69[13]),
    .c(al_591ecc80[6]),
    .o(al_f78b30ce[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c8f379b9 (
    .a(al_2878e2ee),
    .b(al_86280a69[14]),
    .c(al_591ecc80[7]),
    .o(al_f78b30ce[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2414d95e (
    .a(al_2878e2ee),
    .b(al_86280a69[15]),
    .c(al_591ecc80[8]),
    .o(al_f78b30ce[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_54a0fba0 (
    .a(al_2878e2ee),
    .b(al_86280a69[16]),
    .c(al_591ecc80[9]),
    .o(al_f78b30ce[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_54d03012 (
    .a(al_2878e2ee),
    .b(al_86280a69[17]),
    .c(al_591ecc80[10]),
    .o(al_f78b30ce[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f80b2e6b (
    .a(al_2878e2ee),
    .b(al_86280a69[18]),
    .c(al_591ecc80[11]),
    .o(al_f78b30ce[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4287a86b (
    .a(al_2878e2ee),
    .b(al_86280a69[19]),
    .c(al_591ecc80[12]),
    .o(al_f78b30ce[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_62e5b987 (
    .a(al_2878e2ee),
    .b(al_86280a69[20]),
    .c(al_591ecc80[13]),
    .o(al_f78b30ce[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6ce6500e (
    .a(al_2878e2ee),
    .b(al_86280a69[21]),
    .c(al_591ecc80[14]),
    .o(al_f78b30ce[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c8b4913f (
    .a(al_2878e2ee),
    .b(al_86280a69[22]),
    .c(al_591ecc80[15]),
    .o(al_f78b30ce[22]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4cef2c6f (
    .a(al_3029c49a[34]),
    .b(al_3029c49a[35]),
    .c(al_3029c49a[36]),
    .d(al_3029c49a[37]),
    .e(al_3029c49a[38]),
    .f(al_591ecc80[25]),
    .o(al_3a745b61));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_99a53fea (
    .a(al_3a745b61),
    .b(al_3029c49a[32]),
    .c(al_3029c49a[33]),
    .o(al_2878e2ee));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d6da71e (
    .a(al_2878e2ee),
    .b(al_86280a69[23]),
    .c(al_591ecc80[16]),
    .o(al_f78b30ce[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1675244a (
    .a(al_2878e2ee),
    .b(al_86280a69[24]),
    .c(al_591ecc80[17]),
    .o(al_f78b30ce[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_98f73b9d (
    .a(al_2878e2ee),
    .b(al_86280a69[25]),
    .c(al_591ecc80[18]),
    .o(al_f78b30ce[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dca85609 (
    .a(al_2878e2ee),
    .b(al_86280a69[26]),
    .c(al_591ecc80[19]),
    .o(al_f78b30ce[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d67ab856 (
    .a(al_2878e2ee),
    .b(al_86280a69[27]),
    .c(al_591ecc80[20]),
    .o(al_f78b30ce[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_719b035e (
    .a(al_2878e2ee),
    .b(al_86280a69[28]),
    .c(al_591ecc80[21]),
    .o(al_f78b30ce[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e91bee6 (
    .a(al_2878e2ee),
    .b(al_86280a69[29]),
    .c(al_591ecc80[22]),
    .o(al_f78b30ce[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d2e82af9 (
    .a(al_2878e2ee),
    .b(al_86280a69[30]),
    .c(al_591ecc80[23]),
    .o(al_f78b30ce[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e90ef1b (
    .a(al_2878e2ee),
    .b(al_86280a69[31]),
    .c(al_591ecc80[24]),
    .o(al_f78b30ce[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_84f5fce (
    .a(al_2878e2ee),
    .b(al_86280a69[7]),
    .c(al_591ecc80[0]),
    .o(al_f78b30ce[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_892ac0a6 (
    .a(al_2878e2ee),
    .b(al_86280a69[8]),
    .c(al_591ecc80[1]),
    .o(al_f78b30ce[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ba6cdfb9 (
    .a(al_2878e2ee),
    .b(al_86280a69[9]),
    .c(al_591ecc80[2]),
    .o(al_f78b30ce[9]));
  AL_DFF_X al_837001c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0dc7e9e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bade9fae[0]));
  AL_DFF_X al_9cc9fe2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[8]));
  AL_DFF_X al_41b6a3d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[9]));
  AL_DFF_X al_4b5eb6ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[10]));
  AL_DFF_X al_8cc4db69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[11]));
  AL_DFF_X al_3a1606ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[12]));
  AL_DFF_X al_2ff9bbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[13]));
  AL_DFF_X al_14c7ebe8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[14]));
  AL_DFF_X al_ad9101f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[15]));
  AL_DFF_X al_f67ed51d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[16]));
  AL_DFF_X al_743a6b6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[17]));
  AL_DFF_X al_7556b1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[18]));
  AL_DFF_X al_e2254fe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[19]));
  AL_DFF_X al_e5fc68c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[20]));
  AL_DFF_X al_813d0233 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[21]));
  AL_DFF_X al_d56ac716 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[22]));
  AL_DFF_X al_8f89ab02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[23]));
  AL_DFF_X al_9a96c61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[24]));
  AL_DFF_X al_36135b6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[25]));
  AL_DFF_X al_8fb1791b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[26]));
  AL_DFF_X al_d2108ba3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[27]));
  AL_DFF_X al_968a5d74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[28]));
  AL_DFF_X al_e1ea5710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[29]));
  AL_DFF_X al_22a2b910 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[30]));
  AL_DFF_X al_842a5194 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[31]));
  AL_DFF_X al_5a08761d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[32]));
  AL_DFF_X al_20bca572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[33]));
  AL_DFF_X al_ac358971 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[34]));
  AL_DFF_X al_7afe0091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[35]));
  AL_DFF_X al_1d288841 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[36]));
  AL_DFF_X al_8c9ee74a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[37]));
  AL_DFF_X al_c6c5fc3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[6]));
  AL_DFF_X al_58dfc6c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[7]));
  AL_DFF_X al_20229aae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[8]));
  AL_DFF_X al_a4e85ca2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[9]));
  AL_DFF_X al_3b6121ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[10]));
  AL_DFF_X al_5bb8bbec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[11]));
  AL_DFF_X al_a1731e5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[12]));
  AL_DFF_X al_ffe322f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[13]));
  AL_DFF_X al_2a2a6015 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[14]));
  AL_DFF_X al_903c959 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[15]));
  AL_DFF_X al_b35b11c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[16]));
  AL_DFF_X al_e66634a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[17]));
  AL_DFF_X al_734dedd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[0]));
  AL_DFF_X al_1d55b86f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[18]));
  AL_DFF_X al_d2978085 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[19]));
  AL_DFF_X al_a5029241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[20]));
  AL_DFF_X al_3225c616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[21]));
  AL_DFF_X al_1eca4dfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[22]));
  AL_DFF_X al_aaabfc10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[23]));
  AL_DFF_X al_a222ce62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[24]));
  AL_DFF_X al_318e272a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[25]));
  AL_DFF_X al_cdb0a74f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[26]));
  AL_DFF_X al_17b05c47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[27]));
  AL_DFF_X al_e00e97dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[1]));
  AL_DFF_X al_617c9de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[28]));
  AL_DFF_X al_d6b0cc83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[29]));
  AL_DFF_X al_967799ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[30]));
  AL_DFF_X al_85751754 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[31]));
  AL_DFF_X al_ab827abd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[2]));
  AL_DFF_X al_e0383a40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[3]));
  AL_DFF_X al_e11dd453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[4]));
  AL_DFF_X al_1d437ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[5]));
  AL_DFF_X al_1e5e14e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[6]));
  AL_DFF_X al_473fb12d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[7]));
  AL_DFF_X al_13ec4a48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[8]));
  AL_DFF_X al_295e0f37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[9]));
  AL_DFF_X al_6a72b76b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[10]));
  AL_DFF_X al_de98538c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[11]));
  AL_DFF_X al_882f209f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[12]));
  AL_DFF_X al_5f895b8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[13]));
  AL_DFF_X al_2cbbf44d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[14]));
  AL_DFF_X al_bf87e570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[15]));
  AL_DFF_X al_d274328d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[16]));
  AL_DFF_X al_475e97c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[17]));
  AL_DFF_X al_3b5df271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2878e2ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[0]));
  AL_DFF_X al_286fb8e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[18]));
  AL_DFF_X al_12d1f891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[19]));
  AL_DFF_X al_64a1881 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[20]));
  AL_DFF_X al_c26eb920 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[21]));
  AL_DFF_X al_d7cfaa11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[22]));
  AL_DFF_X al_3db4f35f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[23]));
  AL_DFF_X al_e95cdcec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[24]));
  AL_DFF_X al_c754fba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[1]));
  AL_DFF_X al_763d3b41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[2]));
  AL_DFF_X al_1dd0cc13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[3]));
  AL_DFF_X al_b18c22b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[4]));
  AL_DFF_X al_9b97b2cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[5]));
  AL_DFF_X al_318a610e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[6]));
  AL_DFF_X al_65f446fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1431b6e2 (
    .a(1'b0),
    .o({al_1abbaba6,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_34915141 (
    .a(al_9e3033a4[6]),
    .b(al_5181785e[6]),
    .c(al_1abbaba6),
    .o({al_ec19d56e,al_b677b8b1[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce02da5a (
    .a(al_9e3033a4[7]),
    .b(al_5181785e[7]),
    .c(al_ec19d56e),
    .o({al_6409430b,al_b677b8b1[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9e02b10 (
    .a(al_9e3033a4[8]),
    .b(al_5181785e[8]),
    .c(al_6409430b),
    .o({al_33374be5,al_b677b8b1[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_558182ff (
    .a(al_9e3033a4[9]),
    .b(al_5181785e[9]),
    .c(al_33374be5),
    .o({al_97f76d83,al_b677b8b1[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8a8be55 (
    .a(al_9e3033a4[10]),
    .b(al_5181785e[10]),
    .c(al_97f76d83),
    .o({al_111f57ad,al_b677b8b1[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b174c859 (
    .a(al_9e3033a4[11]),
    .b(al_5181785e[11]),
    .c(al_111f57ad),
    .o({al_dd5d3b13,al_b677b8b1[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4fc730f1 (
    .a(al_9e3033a4[12]),
    .b(al_5181785e[12]),
    .c(al_dd5d3b13),
    .o({al_daa9922c,al_b677b8b1[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e81ce80 (
    .a(al_9e3033a4[13]),
    .b(al_5181785e[13]),
    .c(al_daa9922c),
    .o({al_d0a99602,al_b677b8b1[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7dbbe12a (
    .a(al_9e3033a4[14]),
    .b(al_5181785e[14]),
    .c(al_d0a99602),
    .o({al_5a02bf80,al_b677b8b1[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef7f53e5 (
    .a(al_9e3033a4[15]),
    .b(al_5181785e[15]),
    .c(al_5a02bf80),
    .o({al_67d1c21c,al_b677b8b1[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1ca24f0 (
    .a(al_9e3033a4[16]),
    .b(al_5181785e[16]),
    .c(al_67d1c21c),
    .o({al_e79544d1,al_b677b8b1[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5c880745 (
    .a(al_9e3033a4[17]),
    .b(al_5181785e[17]),
    .c(al_e79544d1),
    .o({al_8f3b225e,al_b677b8b1[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be06bc20 (
    .a(al_9e3033a4[18]),
    .b(al_5181785e[18]),
    .c(al_8f3b225e),
    .o({al_b10d3e54,al_b677b8b1[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_643ffb5b (
    .a(al_9e3033a4[19]),
    .b(al_5181785e[19]),
    .c(al_b10d3e54),
    .o({al_fa88be3f,al_b677b8b1[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff8d628b (
    .a(al_9e3033a4[20]),
    .b(al_5181785e[20]),
    .c(al_fa88be3f),
    .o({al_17625a21,al_b677b8b1[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_83dcf7e2 (
    .a(al_9e3033a4[21]),
    .b(al_5181785e[21]),
    .c(al_17625a21),
    .o({al_19e00ab1,al_b677b8b1[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_51b5ea58 (
    .a(al_9e3033a4[22]),
    .b(al_5181785e[22]),
    .c(al_19e00ab1),
    .o({al_c7f6f4df,al_b677b8b1[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f4dfb52 (
    .a(al_9e3033a4[23]),
    .b(al_5181785e[23]),
    .c(al_c7f6f4df),
    .o({al_ea4ffb3c,al_b677b8b1[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_35d964af (
    .a(al_9e3033a4[24]),
    .b(al_5181785e[24]),
    .c(al_ea4ffb3c),
    .o({al_e688eccb,al_b677b8b1[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc1b199f (
    .a(al_9e3033a4[25]),
    .b(al_5181785e[25]),
    .c(al_e688eccb),
    .o({al_ec10f532,al_b677b8b1[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45c76c9e (
    .a(al_9e3033a4[26]),
    .b(al_5181785e[26]),
    .c(al_ec10f532),
    .o({al_a1afdc44,al_b677b8b1[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fafede34 (
    .a(al_9e3033a4[27]),
    .b(al_5181785e[27]),
    .c(al_a1afdc44),
    .o({al_d4e70d9d,al_b677b8b1[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d127216c (
    .a(al_9e3033a4[28]),
    .b(al_5181785e[28]),
    .c(al_d4e70d9d),
    .o({al_16d28d90,al_b677b8b1[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e347c28 (
    .a(al_9e3033a4[29]),
    .b(al_5181785e[29]),
    .c(al_16d28d90),
    .o({al_48808c89,al_b677b8b1[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3db8867 (
    .a(al_9e3033a4[30]),
    .b(al_5181785e[30]),
    .c(al_48808c89),
    .o({al_6216f648,al_b677b8b1[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c439f06 (
    .a(al_9e3033a4[31]),
    .b(al_5181785e[31]),
    .c(al_6216f648),
    .o({al_71a4da9,al_b677b8b1[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_809c0be1 (
    .c(al_71a4da9),
    .o({open_n95,al_b677b8b1[26]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_69d2df8f (
    .a(al_f45fae5e),
    .b(al_9e3033a4[10]),
    .c(al_b677b8b1[4]),
    .o(al_63579c4c[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dc38abb2 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[11]),
    .c(al_b677b8b1[5]),
    .o(al_63579c4c[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_15498e19 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[12]),
    .c(al_b677b8b1[6]),
    .o(al_63579c4c[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfb70fed (
    .a(al_f45fae5e),
    .b(al_9e3033a4[13]),
    .c(al_b677b8b1[7]),
    .o(al_63579c4c[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a22d3c35 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[14]),
    .c(al_b677b8b1[8]),
    .o(al_63579c4c[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5822831f (
    .a(al_f45fae5e),
    .b(al_9e3033a4[15]),
    .c(al_b677b8b1[9]),
    .o(al_63579c4c[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_554930f3 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[16]),
    .c(al_b677b8b1[10]),
    .o(al_63579c4c[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_72a3ff1 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[17]),
    .c(al_b677b8b1[11]),
    .o(al_63579c4c[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9e23b05d (
    .a(al_f45fae5e),
    .b(al_9e3033a4[18]),
    .c(al_b677b8b1[12]),
    .o(al_63579c4c[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_57120ac7 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[19]),
    .c(al_b677b8b1[13]),
    .o(al_63579c4c[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_605e53a1 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[20]),
    .c(al_b677b8b1[14]),
    .o(al_63579c4c[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1e91a57e (
    .a(al_f45fae5e),
    .b(al_9e3033a4[21]),
    .c(al_b677b8b1[15]),
    .o(al_63579c4c[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fd13da36 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[22]),
    .c(al_b677b8b1[16]),
    .o(al_63579c4c[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4e2464d (
    .a(al_f45fae5e),
    .b(al_9e3033a4[23]),
    .c(al_b677b8b1[17]),
    .o(al_63579c4c[23]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_dd9e78f6 (
    .a(al_5181785e[32]),
    .b(al_5181785e[33]),
    .c(al_5181785e[34]),
    .d(al_5181785e[35]),
    .e(al_5181785e[36]),
    .f(al_5181785e[37]),
    .o(al_d7aedbc5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9f8057ca (
    .a(al_d7aedbc5),
    .b(al_b677b8b1[26]),
    .o(al_f45fae5e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_69572de3 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[24]),
    .c(al_b677b8b1[18]),
    .o(al_63579c4c[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e98e59f (
    .a(al_f45fae5e),
    .b(al_9e3033a4[25]),
    .c(al_b677b8b1[19]),
    .o(al_63579c4c[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ef05e4ac (
    .a(al_f45fae5e),
    .b(al_9e3033a4[26]),
    .c(al_b677b8b1[20]),
    .o(al_63579c4c[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7f79dde4 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[27]),
    .c(al_b677b8b1[21]),
    .o(al_63579c4c[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2b64b4b0 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[28]),
    .c(al_b677b8b1[22]),
    .o(al_63579c4c[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1a90d49b (
    .a(al_f45fae5e),
    .b(al_9e3033a4[29]),
    .c(al_b677b8b1[23]),
    .o(al_63579c4c[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e9d85ca (
    .a(al_f45fae5e),
    .b(al_9e3033a4[30]),
    .c(al_b677b8b1[24]),
    .o(al_63579c4c[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bae6af86 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[31]),
    .c(al_b677b8b1[25]),
    .o(al_63579c4c[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_528807c8 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[6]),
    .c(al_b677b8b1[0]),
    .o(al_63579c4c[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5ffaa1a6 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[7]),
    .c(al_b677b8b1[1]),
    .o(al_63579c4c[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5ff7ba0e (
    .a(al_f45fae5e),
    .b(al_9e3033a4[8]),
    .c(al_b677b8b1[2]),
    .o(al_63579c4c[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de82fc64 (
    .a(al_f45fae5e),
    .b(al_9e3033a4[9]),
    .c(al_b677b8b1[3]),
    .o(al_63579c4c[9]));
  AL_DFF_X al_ac39a946 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bade9fae[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f9ab06[0]));
  AL_DFF_X al_7adc28d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[8]));
  AL_DFF_X al_f40ba6f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[9]));
  AL_DFF_X al_e4e13e58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[10]));
  AL_DFF_X al_a658107b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[11]));
  AL_DFF_X al_906782a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[12]));
  AL_DFF_X al_fc6d964 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[13]));
  AL_DFF_X al_2f7ba433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[14]));
  AL_DFF_X al_e60169b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[15]));
  AL_DFF_X al_5531692b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[16]));
  AL_DFF_X al_70a7335c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[17]));
  AL_DFF_X al_1ab01921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[18]));
  AL_DFF_X al_5e02cd78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[19]));
  AL_DFF_X al_4d3c560a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[20]));
  AL_DFF_X al_28177f4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[21]));
  AL_DFF_X al_66d5d441 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[22]));
  AL_DFF_X al_5bb4ee70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[23]));
  AL_DFF_X al_440a5ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[24]));
  AL_DFF_X al_3dd55649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[25]));
  AL_DFF_X al_80b90840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[26]));
  AL_DFF_X al_1f124b8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[27]));
  AL_DFF_X al_ae58e3fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[28]));
  AL_DFF_X al_d54d587d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[29]));
  AL_DFF_X al_aaecde8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[30]));
  AL_DFF_X al_3ecddef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[31]));
  AL_DFF_X al_a45d1d27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[32]));
  AL_DFF_X al_53bbce56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[33]));
  AL_DFF_X al_a7438fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[34]));
  AL_DFF_X al_8bc0403d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[35]));
  AL_DFF_X al_c1065794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[36]));
  AL_DFF_X al_f51320b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[5]));
  AL_DFF_X al_e71fb271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[6]));
  AL_DFF_X al_2b73a0e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[7]));
  AL_DFF_X al_520bb875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[8]));
  AL_DFF_X al_5ef1e75a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[9]));
  AL_DFF_X al_7a4297e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[10]));
  AL_DFF_X al_ea986da7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[11]));
  AL_DFF_X al_74cc8ae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[12]));
  AL_DFF_X al_2d60cd35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[13]));
  AL_DFF_X al_383659d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[14]));
  AL_DFF_X al_7b34e04e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[15]));
  AL_DFF_X al_af640cf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[16]));
  AL_DFF_X al_ec472b93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[17]));
  AL_DFF_X al_c04cfd1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[0]));
  AL_DFF_X al_489c1935 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[18]));
  AL_DFF_X al_3e787941 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[19]));
  AL_DFF_X al_9e64e4f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[20]));
  AL_DFF_X al_b71a0063 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[21]));
  AL_DFF_X al_2fb88ac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[22]));
  AL_DFF_X al_cda30348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[23]));
  AL_DFF_X al_7e4c36b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[24]));
  AL_DFF_X al_8b88f9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[25]));
  AL_DFF_X al_86114405 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[26]));
  AL_DFF_X al_5de5a215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[27]));
  AL_DFF_X al_138cf415 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[1]));
  AL_DFF_X al_c251afb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[28]));
  AL_DFF_X al_8aa4f252 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[29]));
  AL_DFF_X al_7de74184 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[30]));
  AL_DFF_X al_95084e66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[31]));
  AL_DFF_X al_86a1a515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[2]));
  AL_DFF_X al_3f5dfb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[3]));
  AL_DFF_X al_431f965a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[4]));
  AL_DFF_X al_71434deb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[5]));
  AL_DFF_X al_bb43b331 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[6]));
  AL_DFF_X al_95642bf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[7]));
  AL_DFF_X al_f3b684e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[8]));
  AL_DFF_X al_a42247ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[9]));
  AL_DFF_X al_399d1eaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[10]));
  AL_DFF_X al_87213b80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[11]));
  AL_DFF_X al_20e35982 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[12]));
  AL_DFF_X al_6478a9d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[13]));
  AL_DFF_X al_48382f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[14]));
  AL_DFF_X al_d5131777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[15]));
  AL_DFF_X al_69a4ed59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[16]));
  AL_DFF_X al_6d44e6c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[17]));
  AL_DFF_X al_b8e96f4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f45fae5e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[0]));
  AL_DFF_X al_9fbecd47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[18]));
  AL_DFF_X al_d35f5b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[19]));
  AL_DFF_X al_52dcc9d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[20]));
  AL_DFF_X al_982ef376 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[21]));
  AL_DFF_X al_30152ac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[22]));
  AL_DFF_X al_e6505642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[23]));
  AL_DFF_X al_7508b411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[24]));
  AL_DFF_X al_45cfb884 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[25]));
  AL_DFF_X al_a8f3b002 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[1]));
  AL_DFF_X al_910ad0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[2]));
  AL_DFF_X al_da885864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[3]));
  AL_DFF_X al_67cd2ae4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[4]));
  AL_DFF_X al_39e73a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[5]));
  AL_DFF_X al_40f9ddfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[6]));
  AL_DFF_X al_e3ba2ea0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d097171 (
    .a(1'b0),
    .o({al_754bf737,open_n98}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9e2f3300 (
    .a(al_7397600a[5]),
    .b(al_6a56028d[5]),
    .c(al_754bf737),
    .o({al_7fd7f68e,al_64d71d5a[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc730937 (
    .a(al_7397600a[6]),
    .b(al_6a56028d[6]),
    .c(al_7fd7f68e),
    .o({al_b3ed3b7d,al_64d71d5a[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a0b48d96 (
    .a(al_7397600a[7]),
    .b(al_6a56028d[7]),
    .c(al_b3ed3b7d),
    .o({al_c41f5a7c,al_64d71d5a[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_77397675 (
    .a(al_7397600a[8]),
    .b(al_6a56028d[8]),
    .c(al_c41f5a7c),
    .o({al_f31b3480,al_64d71d5a[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14784742 (
    .a(al_7397600a[9]),
    .b(al_6a56028d[9]),
    .c(al_f31b3480),
    .o({al_864bc6dc,al_64d71d5a[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d51f4dd (
    .a(al_7397600a[10]),
    .b(al_6a56028d[10]),
    .c(al_864bc6dc),
    .o({al_f693e61d,al_64d71d5a[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f723467 (
    .a(al_7397600a[11]),
    .b(al_6a56028d[11]),
    .c(al_f693e61d),
    .o({al_47955db6,al_64d71d5a[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2e2500 (
    .a(al_7397600a[12]),
    .b(al_6a56028d[12]),
    .c(al_47955db6),
    .o({al_cc078df4,al_64d71d5a[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5aa1d15a (
    .a(al_7397600a[13]),
    .b(al_6a56028d[13]),
    .c(al_cc078df4),
    .o({al_58dab36d,al_64d71d5a[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_698c457e (
    .a(al_7397600a[14]),
    .b(al_6a56028d[14]),
    .c(al_58dab36d),
    .o({al_3e035452,al_64d71d5a[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cef124b5 (
    .a(al_7397600a[15]),
    .b(al_6a56028d[15]),
    .c(al_3e035452),
    .o({al_106a827,al_64d71d5a[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f130734c (
    .a(al_7397600a[16]),
    .b(al_6a56028d[16]),
    .c(al_106a827),
    .o({al_f709c5ab,al_64d71d5a[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_330b2e33 (
    .a(al_7397600a[17]),
    .b(al_6a56028d[17]),
    .c(al_f709c5ab),
    .o({al_56abe384,al_64d71d5a[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6230e8f2 (
    .a(al_7397600a[18]),
    .b(al_6a56028d[18]),
    .c(al_56abe384),
    .o({al_7418c94f,al_64d71d5a[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d2812258 (
    .a(al_7397600a[19]),
    .b(al_6a56028d[19]),
    .c(al_7418c94f),
    .o({al_efa49dac,al_64d71d5a[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b9d7159e (
    .a(al_7397600a[20]),
    .b(al_6a56028d[20]),
    .c(al_efa49dac),
    .o({al_e130ad23,al_64d71d5a[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1bd3436f (
    .a(al_7397600a[21]),
    .b(al_6a56028d[21]),
    .c(al_e130ad23),
    .o({al_2f299606,al_64d71d5a[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5d133bf (
    .a(al_7397600a[22]),
    .b(al_6a56028d[22]),
    .c(al_2f299606),
    .o({al_925eb901,al_64d71d5a[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8c659c63 (
    .a(al_7397600a[23]),
    .b(al_6a56028d[23]),
    .c(al_925eb901),
    .o({al_daeef93a,al_64d71d5a[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33f675fd (
    .a(al_7397600a[24]),
    .b(al_6a56028d[24]),
    .c(al_daeef93a),
    .o({al_2ff932f4,al_64d71d5a[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7551e068 (
    .a(al_7397600a[25]),
    .b(al_6a56028d[25]),
    .c(al_2ff932f4),
    .o({al_2e6e4c5b,al_64d71d5a[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_11eb7df7 (
    .a(al_7397600a[26]),
    .b(al_6a56028d[26]),
    .c(al_2e6e4c5b),
    .o({al_2a6886e2,al_64d71d5a[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4549d1d3 (
    .a(al_7397600a[27]),
    .b(al_6a56028d[27]),
    .c(al_2a6886e2),
    .o({al_1f220fb,al_64d71d5a[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c3678be (
    .a(al_7397600a[28]),
    .b(al_6a56028d[28]),
    .c(al_1f220fb),
    .o({al_7154b9a7,al_64d71d5a[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47a8dbd1 (
    .a(al_7397600a[29]),
    .b(al_6a56028d[29]),
    .c(al_7154b9a7),
    .o({al_1bf81a9b,al_64d71d5a[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_77a2169e (
    .a(al_7397600a[30]),
    .b(al_6a56028d[30]),
    .c(al_1bf81a9b),
    .o({al_1b451831,al_64d71d5a[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d2b6579a (
    .a(al_7397600a[31]),
    .b(al_6a56028d[31]),
    .c(al_1b451831),
    .o({al_72e17b7c,al_64d71d5a[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_948e069b (
    .c(al_72e17b7c),
    .o({open_n101,al_64d71d5a[27]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5c5d1279 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[10]),
    .c(al_64d71d5a[5]),
    .o(al_2c297489[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a1399fe8 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[11]),
    .c(al_64d71d5a[6]),
    .o(al_2c297489[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ddc6f7f7 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[12]),
    .c(al_64d71d5a[7]),
    .o(al_2c297489[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_77c334a (
    .a(al_a1fc4ea8),
    .b(al_7397600a[13]),
    .c(al_64d71d5a[8]),
    .o(al_2c297489[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d3add3dd (
    .a(al_a1fc4ea8),
    .b(al_7397600a[14]),
    .c(al_64d71d5a[9]),
    .o(al_2c297489[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e7d9867 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[15]),
    .c(al_64d71d5a[10]),
    .o(al_2c297489[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e78b10e (
    .a(al_a1fc4ea8),
    .b(al_7397600a[16]),
    .c(al_64d71d5a[11]),
    .o(al_2c297489[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e740a918 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[17]),
    .c(al_64d71d5a[12]),
    .o(al_2c297489[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99bfcbf4 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[18]),
    .c(al_64d71d5a[13]),
    .o(al_2c297489[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1d06849e (
    .a(al_a1fc4ea8),
    .b(al_7397600a[19]),
    .c(al_64d71d5a[14]),
    .o(al_2c297489[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_88021601 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[20]),
    .c(al_64d71d5a[15]),
    .o(al_2c297489[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_285f8831 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[21]),
    .c(al_64d71d5a[16]),
    .o(al_2c297489[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6034d936 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[22]),
    .c(al_64d71d5a[17]),
    .o(al_2c297489[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f11b9504 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[23]),
    .c(al_64d71d5a[18]),
    .o(al_2c297489[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e50e5e88 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[24]),
    .c(al_64d71d5a[19]),
    .o(al_2c297489[24]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_948dbf8d (
    .a(al_6a56028d[32]),
    .b(al_6a56028d[33]),
    .c(al_6a56028d[34]),
    .d(al_6a56028d[35]),
    .e(al_6a56028d[36]),
    .f(al_64d71d5a[27]),
    .o(al_a1fc4ea8));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3c29dfb4 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[25]),
    .c(al_64d71d5a[20]),
    .o(al_2c297489[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_be4fad80 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[26]),
    .c(al_64d71d5a[21]),
    .o(al_2c297489[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d88731a4 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[27]),
    .c(al_64d71d5a[22]),
    .o(al_2c297489[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2a8943 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[28]),
    .c(al_64d71d5a[23]),
    .o(al_2c297489[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a1786b68 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[29]),
    .c(al_64d71d5a[24]),
    .o(al_2c297489[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93f2f040 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[30]),
    .c(al_64d71d5a[25]),
    .o(al_2c297489[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_84afee8 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[31]),
    .c(al_64d71d5a[26]),
    .o(al_2c297489[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d2f59bf1 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[5]),
    .c(al_64d71d5a[0]),
    .o(al_2c297489[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a24a0bf4 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[6]),
    .c(al_64d71d5a[1]),
    .o(al_2c297489[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b22a21be (
    .a(al_a1fc4ea8),
    .b(al_7397600a[7]),
    .c(al_64d71d5a[2]),
    .o(al_2c297489[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e67b0a4f (
    .a(al_a1fc4ea8),
    .b(al_7397600a[8]),
    .c(al_64d71d5a[3]),
    .o(al_2c297489[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a982d554 (
    .a(al_a1fc4ea8),
    .b(al_7397600a[9]),
    .c(al_64d71d5a[4]),
    .o(al_2c297489[9]));
  AL_DFF_X al_a01bdf6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8f9ab06[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fee4bd37[0]));
  AL_DFF_X al_357f1a32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[8]));
  AL_DFF_X al_9a776ea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[9]));
  AL_DFF_X al_b0e4fd80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[10]));
  AL_DFF_X al_cc3f7e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[11]));
  AL_DFF_X al_8da5e71e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[12]));
  AL_DFF_X al_61afd285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[13]));
  AL_DFF_X al_94f89e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[14]));
  AL_DFF_X al_d811b449 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[15]));
  AL_DFF_X al_ed9b689f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[16]));
  AL_DFF_X al_8e8cdbaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[17]));
  AL_DFF_X al_b338e1d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[18]));
  AL_DFF_X al_24867b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[19]));
  AL_DFF_X al_155b5c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[20]));
  AL_DFF_X al_40a55559 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[21]));
  AL_DFF_X al_a8cb326d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[22]));
  AL_DFF_X al_56f0bd9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[23]));
  AL_DFF_X al_3dc2501e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[24]));
  AL_DFF_X al_e067fd4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[25]));
  AL_DFF_X al_658489ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[26]));
  AL_DFF_X al_4d4743c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[27]));
  AL_DFF_X al_d287c6f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[28]));
  AL_DFF_X al_2330cbb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[29]));
  AL_DFF_X al_44e25ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[30]));
  AL_DFF_X al_73411bd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[31]));
  AL_DFF_X al_508049fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[32]));
  AL_DFF_X al_9d67371e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[33]));
  AL_DFF_X al_34b61ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[34]));
  AL_DFF_X al_5a19486e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[35]));
  AL_DFF_X al_4a779f04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[4]));
  AL_DFF_X al_aea4d16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[5]));
  AL_DFF_X al_57c3d7dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[6]));
  AL_DFF_X al_5092fed6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[7]));
  AL_DFF_X al_ff50b69e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[8]));
  AL_DFF_X al_542c5466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[9]));
  AL_DFF_X al_d711901b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[10]));
  AL_DFF_X al_fb38d079 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[11]));
  AL_DFF_X al_606807 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[12]));
  AL_DFF_X al_34b40683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[13]));
  AL_DFF_X al_85e05024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[14]));
  AL_DFF_X al_e942dcff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[15]));
  AL_DFF_X al_dc0c05a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[16]));
  AL_DFF_X al_c656a86f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[17]));
  AL_DFF_X al_b51d9aa4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[0]));
  AL_DFF_X al_6834f9fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[18]));
  AL_DFF_X al_ec83082b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[19]));
  AL_DFF_X al_3db9e412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[20]));
  AL_DFF_X al_899cbb99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[21]));
  AL_DFF_X al_71379287 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[22]));
  AL_DFF_X al_c6605c29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[23]));
  AL_DFF_X al_91152122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[24]));
  AL_DFF_X al_1bfdc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[25]));
  AL_DFF_X al_3b513970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[26]));
  AL_DFF_X al_d8c1c9d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[27]));
  AL_DFF_X al_e5dd8a9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[1]));
  AL_DFF_X al_a76f7657 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[28]));
  AL_DFF_X al_f2760a29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[29]));
  AL_DFF_X al_313f802b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[30]));
  AL_DFF_X al_cfdb03de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[31]));
  AL_DFF_X al_a5b658e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[2]));
  AL_DFF_X al_d44ccb4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[3]));
  AL_DFF_X al_a8857375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[4]));
  AL_DFF_X al_a3073509 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[5]));
  AL_DFF_X al_7f4d584 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[6]));
  AL_DFF_X al_430193b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[7]));
  AL_DFF_X al_e5afa724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[8]));
  AL_DFF_X al_d5636866 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[9]));
  AL_DFF_X al_c0d76e5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[10]));
  AL_DFF_X al_7b7dc4dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[11]));
  AL_DFF_X al_5ad8e11b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[12]));
  AL_DFF_X al_de7b1d72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[13]));
  AL_DFF_X al_efc4eda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[14]));
  AL_DFF_X al_ede43bde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[15]));
  AL_DFF_X al_e171fd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[16]));
  AL_DFF_X al_c795c975 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[17]));
  AL_DFF_X al_24442eeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a1fc4ea8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[0]));
  AL_DFF_X al_4be4fc87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[18]));
  AL_DFF_X al_f9bda6b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[19]));
  AL_DFF_X al_6357a0d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[20]));
  AL_DFF_X al_1dc8e7f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[21]));
  AL_DFF_X al_ecc97e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[22]));
  AL_DFF_X al_9bd57b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[23]));
  AL_DFF_X al_b1e64020 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[24]));
  AL_DFF_X al_4c27f563 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[25]));
  AL_DFF_X al_d13fa94a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[26]));
  AL_DFF_X al_c4a33bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[1]));
  AL_DFF_X al_d5161d1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[2]));
  AL_DFF_X al_139cf0c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[3]));
  AL_DFF_X al_ea572dee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[4]));
  AL_DFF_X al_94240d41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[5]));
  AL_DFF_X al_4c96883f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[6]));
  AL_DFF_X al_831353ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_97fe3c3a (
    .a(1'b0),
    .o({al_dde82c43,open_n104}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fbb007d9 (
    .a(al_e4be4089[4]),
    .b(al_b6768e55[4]),
    .c(al_dde82c43),
    .o({al_b1d329d9,al_c20bde66[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_71b4340c (
    .a(al_e4be4089[5]),
    .b(al_b6768e55[5]),
    .c(al_b1d329d9),
    .o({al_c8aee28f,al_c20bde66[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_445114cd (
    .a(al_e4be4089[6]),
    .b(al_b6768e55[6]),
    .c(al_c8aee28f),
    .o({al_b33e7544,al_c20bde66[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_807224fc (
    .a(al_e4be4089[7]),
    .b(al_b6768e55[7]),
    .c(al_b33e7544),
    .o({al_accca793,al_c20bde66[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_87a4e3fd (
    .a(al_e4be4089[8]),
    .b(al_b6768e55[8]),
    .c(al_accca793),
    .o({al_4dd25e15,al_c20bde66[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92db03af (
    .a(al_e4be4089[9]),
    .b(al_b6768e55[9]),
    .c(al_4dd25e15),
    .o({al_c76b4c37,al_c20bde66[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1196df5 (
    .a(al_e4be4089[10]),
    .b(al_b6768e55[10]),
    .c(al_c76b4c37),
    .o({al_b7a54e24,al_c20bde66[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ca2df25 (
    .a(al_e4be4089[11]),
    .b(al_b6768e55[11]),
    .c(al_b7a54e24),
    .o({al_85587067,al_c20bde66[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e88365f (
    .a(al_e4be4089[12]),
    .b(al_b6768e55[12]),
    .c(al_85587067),
    .o({al_1ff06f87,al_c20bde66[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9fc9481c (
    .a(al_e4be4089[13]),
    .b(al_b6768e55[13]),
    .c(al_1ff06f87),
    .o({al_143fe859,al_c20bde66[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6c471e48 (
    .a(al_e4be4089[14]),
    .b(al_b6768e55[14]),
    .c(al_143fe859),
    .o({al_cd6d2794,al_c20bde66[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_388f0223 (
    .a(al_e4be4089[15]),
    .b(al_b6768e55[15]),
    .c(al_cd6d2794),
    .o({al_e59fc5bd,al_c20bde66[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_46217ab9 (
    .a(al_e4be4089[16]),
    .b(al_b6768e55[16]),
    .c(al_e59fc5bd),
    .o({al_bd4c5933,al_c20bde66[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_77cc2d68 (
    .a(al_e4be4089[17]),
    .b(al_b6768e55[17]),
    .c(al_bd4c5933),
    .o({al_6c260918,al_c20bde66[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e44aa20c (
    .a(al_e4be4089[18]),
    .b(al_b6768e55[18]),
    .c(al_6c260918),
    .o({al_6b532b61,al_c20bde66[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_806c985a (
    .a(al_e4be4089[19]),
    .b(al_b6768e55[19]),
    .c(al_6b532b61),
    .o({al_9cdbacea,al_c20bde66[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e9ebef51 (
    .a(al_e4be4089[20]),
    .b(al_b6768e55[20]),
    .c(al_9cdbacea),
    .o({al_232548,al_c20bde66[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8684231 (
    .a(al_e4be4089[21]),
    .b(al_b6768e55[21]),
    .c(al_232548),
    .o({al_e1d75325,al_c20bde66[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_94ac0fa3 (
    .a(al_e4be4089[22]),
    .b(al_b6768e55[22]),
    .c(al_e1d75325),
    .o({al_87178f5,al_c20bde66[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_24dac0b7 (
    .a(al_e4be4089[23]),
    .b(al_b6768e55[23]),
    .c(al_87178f5),
    .o({al_70012e88,al_c20bde66[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f1a5a6a1 (
    .a(al_e4be4089[24]),
    .b(al_b6768e55[24]),
    .c(al_70012e88),
    .o({al_452820cd,al_c20bde66[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2caa1a5d (
    .a(al_e4be4089[25]),
    .b(al_b6768e55[25]),
    .c(al_452820cd),
    .o({al_392bc465,al_c20bde66[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3b219ec (
    .a(al_e4be4089[26]),
    .b(al_b6768e55[26]),
    .c(al_392bc465),
    .o({al_adc3cec6,al_c20bde66[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c3e4e703 (
    .a(al_e4be4089[27]),
    .b(al_b6768e55[27]),
    .c(al_adc3cec6),
    .o({al_852fa027,al_c20bde66[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e08e8fdd (
    .a(al_e4be4089[28]),
    .b(al_b6768e55[28]),
    .c(al_852fa027),
    .o({al_3c9f5595,al_c20bde66[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a17a283 (
    .a(al_e4be4089[29]),
    .b(al_b6768e55[29]),
    .c(al_3c9f5595),
    .o({al_829de986,al_c20bde66[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50c8448c (
    .a(al_e4be4089[30]),
    .b(al_b6768e55[30]),
    .c(al_829de986),
    .o({al_e3bf1d53,al_c20bde66[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_20beb8fe (
    .a(al_e4be4089[31]),
    .b(al_b6768e55[31]),
    .c(al_e3bf1d53),
    .o({al_e6964d98,al_c20bde66[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e240eb9 (
    .c(al_e6964d98),
    .o({open_n107,al_c20bde66[28]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8c6d1bd5 (
    .a(al_188e472a),
    .b(al_e4be4089[10]),
    .c(al_c20bde66[6]),
    .o(al_9857f6b5[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_afc05270 (
    .a(al_188e472a),
    .b(al_e4be4089[11]),
    .c(al_c20bde66[7]),
    .o(al_9857f6b5[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dbf784a1 (
    .a(al_188e472a),
    .b(al_e4be4089[12]),
    .c(al_c20bde66[8]),
    .o(al_9857f6b5[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e3bfc2a0 (
    .a(al_188e472a),
    .b(al_e4be4089[13]),
    .c(al_c20bde66[9]),
    .o(al_9857f6b5[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_94e8ff88 (
    .a(al_188e472a),
    .b(al_e4be4089[14]),
    .c(al_c20bde66[10]),
    .o(al_9857f6b5[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ca38a50 (
    .a(al_188e472a),
    .b(al_e4be4089[15]),
    .c(al_c20bde66[11]),
    .o(al_9857f6b5[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a21b20e7 (
    .a(al_188e472a),
    .b(al_e4be4089[16]),
    .c(al_c20bde66[12]),
    .o(al_9857f6b5[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_13959bb1 (
    .a(al_188e472a),
    .b(al_e4be4089[17]),
    .c(al_c20bde66[13]),
    .o(al_9857f6b5[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_10ceec37 (
    .a(al_188e472a),
    .b(al_e4be4089[18]),
    .c(al_c20bde66[14]),
    .o(al_9857f6b5[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4cb4e9fc (
    .a(al_188e472a),
    .b(al_e4be4089[19]),
    .c(al_c20bde66[15]),
    .o(al_9857f6b5[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_812d1ca8 (
    .a(al_188e472a),
    .b(al_e4be4089[20]),
    .c(al_c20bde66[16]),
    .o(al_9857f6b5[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ce868b8d (
    .a(al_188e472a),
    .b(al_e4be4089[21]),
    .c(al_c20bde66[17]),
    .o(al_9857f6b5[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34b7cb0f (
    .a(al_188e472a),
    .b(al_e4be4089[22]),
    .c(al_c20bde66[18]),
    .o(al_9857f6b5[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aeb1fe37 (
    .a(al_188e472a),
    .b(al_e4be4089[23]),
    .c(al_c20bde66[19]),
    .o(al_9857f6b5[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_162fda05 (
    .a(al_188e472a),
    .b(al_e4be4089[24]),
    .c(al_c20bde66[20]),
    .o(al_9857f6b5[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0639d5d (
    .a(al_188e472a),
    .b(al_e4be4089[25]),
    .c(al_c20bde66[21]),
    .o(al_9857f6b5[25]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_255f48b6 (
    .a(al_b6768e55[32]),
    .b(al_b6768e55[33]),
    .c(al_b6768e55[34]),
    .d(al_b6768e55[35]),
    .e(al_c20bde66[28]),
    .o(al_188e472a));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ce09416f (
    .a(al_188e472a),
    .b(al_e4be4089[26]),
    .c(al_c20bde66[22]),
    .o(al_9857f6b5[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dd419afc (
    .a(al_188e472a),
    .b(al_e4be4089[27]),
    .c(al_c20bde66[23]),
    .o(al_9857f6b5[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2f3c91a (
    .a(al_188e472a),
    .b(al_e4be4089[28]),
    .c(al_c20bde66[24]),
    .o(al_9857f6b5[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_601e8e7a (
    .a(al_188e472a),
    .b(al_e4be4089[29]),
    .c(al_c20bde66[25]),
    .o(al_9857f6b5[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7ac0d4fa (
    .a(al_188e472a),
    .b(al_e4be4089[30]),
    .c(al_c20bde66[26]),
    .o(al_9857f6b5[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_65aa7b93 (
    .a(al_188e472a),
    .b(al_e4be4089[31]),
    .c(al_c20bde66[27]),
    .o(al_9857f6b5[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee4d2a90 (
    .a(al_188e472a),
    .b(al_e4be4089[4]),
    .c(al_c20bde66[0]),
    .o(al_9857f6b5[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_66a90317 (
    .a(al_188e472a),
    .b(al_e4be4089[5]),
    .c(al_c20bde66[1]),
    .o(al_9857f6b5[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f2cd2814 (
    .a(al_188e472a),
    .b(al_e4be4089[6]),
    .c(al_c20bde66[2]),
    .o(al_9857f6b5[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c7cf0834 (
    .a(al_188e472a),
    .b(al_e4be4089[7]),
    .c(al_c20bde66[3]),
    .o(al_9857f6b5[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a31e4289 (
    .a(al_188e472a),
    .b(al_e4be4089[8]),
    .c(al_c20bde66[4]),
    .o(al_9857f6b5[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7422d80 (
    .a(al_188e472a),
    .b(al_e4be4089[9]),
    .c(al_c20bde66[5]),
    .o(al_9857f6b5[9]));
  AL_DFF_X al_db9ef6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fee4bd37[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e0e2aae4[0]));
  AL_DFF_X al_744243ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[8]));
  AL_DFF_X al_b3609633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[9]));
  AL_DFF_X al_7a8867fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[10]));
  AL_DFF_X al_3fea02c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[11]));
  AL_DFF_X al_557092d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[12]));
  AL_DFF_X al_f3efe660 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[13]));
  AL_DFF_X al_32c90653 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[14]));
  AL_DFF_X al_16c76650 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[15]));
  AL_DFF_X al_d7d7e859 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[16]));
  AL_DFF_X al_306f7c38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[17]));
  AL_DFF_X al_214a1cd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[18]));
  AL_DFF_X al_c4518989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[19]));
  AL_DFF_X al_131f21f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[20]));
  AL_DFF_X al_4e674112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[21]));
  AL_DFF_X al_5c1af8da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[22]));
  AL_DFF_X al_83363eab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[23]));
  AL_DFF_X al_18c36b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[24]));
  AL_DFF_X al_32491724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[25]));
  AL_DFF_X al_b8e07d6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[26]));
  AL_DFF_X al_466a66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[27]));
  AL_DFF_X al_568e3781 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[28]));
  AL_DFF_X al_1748a8f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[29]));
  AL_DFF_X al_52498111 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[30]));
  AL_DFF_X al_93d0de9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[31]));
  AL_DFF_X al_9b80b2f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[32]));
  AL_DFF_X al_19b79172 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[33]));
  AL_DFF_X al_48e1ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[34]));
  AL_DFF_X al_8cd9cf2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[3]));
  AL_DFF_X al_8812fb51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[4]));
  AL_DFF_X al_20ea267a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[5]));
  AL_DFF_X al_a51de33f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[6]));
  AL_DFF_X al_161efd03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[7]));
  AL_DFF_X al_7778ee00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[8]));
  AL_DFF_X al_1a55efc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[9]));
  AL_DFF_X al_3e13bd48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[10]));
  AL_DFF_X al_5bde5b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[11]));
  AL_DFF_X al_2ffb2115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[12]));
  AL_DFF_X al_ba51121f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[13]));
  AL_DFF_X al_5afa016f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[14]));
  AL_DFF_X al_4bfd5a26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[15]));
  AL_DFF_X al_f78cc6dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[16]));
  AL_DFF_X al_913239f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[17]));
  AL_DFF_X al_82ce4c19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[0]));
  AL_DFF_X al_d4094e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[18]));
  AL_DFF_X al_322b4f04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[19]));
  AL_DFF_X al_e336a39b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[20]));
  AL_DFF_X al_17e0341e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[21]));
  AL_DFF_X al_b8071361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[22]));
  AL_DFF_X al_3f76117a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[23]));
  AL_DFF_X al_cb97ab5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[24]));
  AL_DFF_X al_49cf54fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[25]));
  AL_DFF_X al_2ba448e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[26]));
  AL_DFF_X al_37e68a19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[27]));
  AL_DFF_X al_ea479ee3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[1]));
  AL_DFF_X al_da38eb6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[28]));
  AL_DFF_X al_8d981788 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[29]));
  AL_DFF_X al_43d41971 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[30]));
  AL_DFF_X al_b6a85e6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[31]));
  AL_DFF_X al_efb4135c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[2]));
  AL_DFF_X al_ff4eb381 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[3]));
  AL_DFF_X al_d5810c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[4]));
  AL_DFF_X al_a059413f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[5]));
  AL_DFF_X al_15dea8ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[6]));
  AL_DFF_X al_507f24c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[7]));
  AL_DFF_X al_314c199e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[8]));
  AL_DFF_X al_4985edbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[9]));
  AL_DFF_X al_61b309d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[10]));
  AL_DFF_X al_f9d32b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[11]));
  AL_DFF_X al_129510d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[12]));
  AL_DFF_X al_17ca42b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[13]));
  AL_DFF_X al_6e33643b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[14]));
  AL_DFF_X al_31a08202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[15]));
  AL_DFF_X al_7c17021f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[16]));
  AL_DFF_X al_dbe14f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[17]));
  AL_DFF_X al_6333d411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_188e472a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[0]));
  AL_DFF_X al_82a0034b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[18]));
  AL_DFF_X al_6dda13d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[19]));
  AL_DFF_X al_fbb5bf43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[20]));
  AL_DFF_X al_d3122d3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[21]));
  AL_DFF_X al_f937dbdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[22]));
  AL_DFF_X al_fd04a76a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[23]));
  AL_DFF_X al_b732b427 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[24]));
  AL_DFF_X al_40fcc083 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[25]));
  AL_DFF_X al_a94b0edc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[26]));
  AL_DFF_X al_abf7920f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[27]));
  AL_DFF_X al_1462305b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[1]));
  AL_DFF_X al_df25482e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[2]));
  AL_DFF_X al_a13909bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[3]));
  AL_DFF_X al_545f9c29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[4]));
  AL_DFF_X al_ccd9624 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[5]));
  AL_DFF_X al_6c9293a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[6]));
  AL_DFF_X al_662a09ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d8358717 (
    .a(1'b0),
    .o({al_d8b8a6e2,open_n110}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9a9a553 (
    .a(al_4a463b38[3]),
    .b(al_222a5f4d[3]),
    .c(al_d8b8a6e2),
    .o({al_8044404c,al_632b75dc[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21c6b0be (
    .a(al_4a463b38[4]),
    .b(al_222a5f4d[4]),
    .c(al_8044404c),
    .o({al_ca8e61e8,al_632b75dc[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e9797f0 (
    .a(al_4a463b38[5]),
    .b(al_222a5f4d[5]),
    .c(al_ca8e61e8),
    .o({al_3144b627,al_632b75dc[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d0a796f (
    .a(al_4a463b38[6]),
    .b(al_222a5f4d[6]),
    .c(al_3144b627),
    .o({al_cb5d4eb2,al_632b75dc[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c73b4123 (
    .a(al_4a463b38[7]),
    .b(al_222a5f4d[7]),
    .c(al_cb5d4eb2),
    .o({al_e2af005f,al_632b75dc[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ecce2016 (
    .a(al_4a463b38[8]),
    .b(al_222a5f4d[8]),
    .c(al_e2af005f),
    .o({al_dd8f16d1,al_632b75dc[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97358cac (
    .a(al_4a463b38[9]),
    .b(al_222a5f4d[9]),
    .c(al_dd8f16d1),
    .o({al_f2a22ed1,al_632b75dc[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b74c802 (
    .a(al_4a463b38[10]),
    .b(al_222a5f4d[10]),
    .c(al_f2a22ed1),
    .o({al_d1a88ad2,al_632b75dc[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aeb99b20 (
    .a(al_4a463b38[11]),
    .b(al_222a5f4d[11]),
    .c(al_d1a88ad2),
    .o({al_3c316ef,al_632b75dc[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b07d80fb (
    .a(al_4a463b38[12]),
    .b(al_222a5f4d[12]),
    .c(al_3c316ef),
    .o({al_a2fff3ec,al_632b75dc[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8a1b838 (
    .a(al_4a463b38[13]),
    .b(al_222a5f4d[13]),
    .c(al_a2fff3ec),
    .o({al_f6ffe199,al_632b75dc[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_683538d4 (
    .a(al_4a463b38[14]),
    .b(al_222a5f4d[14]),
    .c(al_f6ffe199),
    .o({al_aa4c6187,al_632b75dc[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_826988fd (
    .a(al_4a463b38[15]),
    .b(al_222a5f4d[15]),
    .c(al_aa4c6187),
    .o({al_3d105014,al_632b75dc[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f95e76e0 (
    .a(al_4a463b38[16]),
    .b(al_222a5f4d[16]),
    .c(al_3d105014),
    .o({al_f0daa0db,al_632b75dc[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ffd993ac (
    .a(al_4a463b38[17]),
    .b(al_222a5f4d[17]),
    .c(al_f0daa0db),
    .o({al_47c0210d,al_632b75dc[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_656faafe (
    .a(al_4a463b38[18]),
    .b(al_222a5f4d[18]),
    .c(al_47c0210d),
    .o({al_85b1bb55,al_632b75dc[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9cd69d08 (
    .a(al_4a463b38[19]),
    .b(al_222a5f4d[19]),
    .c(al_85b1bb55),
    .o({al_ebd1e7fe,al_632b75dc[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_75f21671 (
    .a(al_4a463b38[20]),
    .b(al_222a5f4d[20]),
    .c(al_ebd1e7fe),
    .o({al_bc14fb86,al_632b75dc[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee8ac2d1 (
    .a(al_4a463b38[21]),
    .b(al_222a5f4d[21]),
    .c(al_bc14fb86),
    .o({al_dd5db619,al_632b75dc[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3a07367 (
    .a(al_4a463b38[22]),
    .b(al_222a5f4d[22]),
    .c(al_dd5db619),
    .o({al_3e3b2341,al_632b75dc[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dbd673f (
    .a(al_4a463b38[23]),
    .b(al_222a5f4d[23]),
    .c(al_3e3b2341),
    .o({al_9b3654ad,al_632b75dc[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6fac8d0 (
    .a(al_4a463b38[24]),
    .b(al_222a5f4d[24]),
    .c(al_9b3654ad),
    .o({al_100303d6,al_632b75dc[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_375191a7 (
    .a(al_4a463b38[25]),
    .b(al_222a5f4d[25]),
    .c(al_100303d6),
    .o({al_50e17485,al_632b75dc[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3cfcf4a7 (
    .a(al_4a463b38[26]),
    .b(al_222a5f4d[26]),
    .c(al_50e17485),
    .o({al_3b8d6cb9,al_632b75dc[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af74aba3 (
    .a(al_4a463b38[27]),
    .b(al_222a5f4d[27]),
    .c(al_3b8d6cb9),
    .o({al_83167981,al_632b75dc[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_faef6e85 (
    .a(al_4a463b38[28]),
    .b(al_222a5f4d[28]),
    .c(al_83167981),
    .o({al_3fb5c0bf,al_632b75dc[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fd867ae (
    .a(al_4a463b38[29]),
    .b(al_222a5f4d[29]),
    .c(al_3fb5c0bf),
    .o({al_f7a0a5e,al_632b75dc[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_849de08c (
    .a(al_4a463b38[30]),
    .b(al_222a5f4d[30]),
    .c(al_f7a0a5e),
    .o({al_28c3840c,al_632b75dc[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f60ba96f (
    .a(al_4a463b38[31]),
    .b(al_222a5f4d[31]),
    .c(al_28c3840c),
    .o({al_a5df252b,al_632b75dc[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_29fe7e80 (
    .c(al_a5df252b),
    .o({open_n113,al_632b75dc[29]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_361b4e1c (
    .a(al_855effe8),
    .b(al_4a463b38[10]),
    .c(al_632b75dc[7]),
    .o(al_e343d659[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cc07d950 (
    .a(al_855effe8),
    .b(al_4a463b38[11]),
    .c(al_632b75dc[8]),
    .o(al_e343d659[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e1c8930a (
    .a(al_855effe8),
    .b(al_4a463b38[12]),
    .c(al_632b75dc[9]),
    .o(al_e343d659[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f2d19280 (
    .a(al_855effe8),
    .b(al_4a463b38[13]),
    .c(al_632b75dc[10]),
    .o(al_e343d659[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_954d45fb (
    .a(al_855effe8),
    .b(al_4a463b38[14]),
    .c(al_632b75dc[11]),
    .o(al_e343d659[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4e2dfab9 (
    .a(al_855effe8),
    .b(al_4a463b38[15]),
    .c(al_632b75dc[12]),
    .o(al_e343d659[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e9b75cc5 (
    .a(al_855effe8),
    .b(al_4a463b38[16]),
    .c(al_632b75dc[13]),
    .o(al_e343d659[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1318a70b (
    .a(al_855effe8),
    .b(al_4a463b38[17]),
    .c(al_632b75dc[14]),
    .o(al_e343d659[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1cfb913b (
    .a(al_855effe8),
    .b(al_4a463b38[18]),
    .c(al_632b75dc[15]),
    .o(al_e343d659[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a97a84a2 (
    .a(al_855effe8),
    .b(al_4a463b38[19]),
    .c(al_632b75dc[16]),
    .o(al_e343d659[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9bc6d77a (
    .a(al_855effe8),
    .b(al_4a463b38[20]),
    .c(al_632b75dc[17]),
    .o(al_e343d659[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4fa5015c (
    .a(al_855effe8),
    .b(al_4a463b38[21]),
    .c(al_632b75dc[18]),
    .o(al_e343d659[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9447a0dd (
    .a(al_855effe8),
    .b(al_4a463b38[22]),
    .c(al_632b75dc[19]),
    .o(al_e343d659[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2cc9bd8 (
    .a(al_855effe8),
    .b(al_4a463b38[23]),
    .c(al_632b75dc[20]),
    .o(al_e343d659[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b7b6b52 (
    .a(al_855effe8),
    .b(al_4a463b38[24]),
    .c(al_632b75dc[21]),
    .o(al_e343d659[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_67fe5ba4 (
    .a(al_855effe8),
    .b(al_4a463b38[25]),
    .c(al_632b75dc[22]),
    .o(al_e343d659[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1fa28c08 (
    .a(al_855effe8),
    .b(al_4a463b38[26]),
    .c(al_632b75dc[23]),
    .o(al_e343d659[26]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8da17227 (
    .a(al_222a5f4d[32]),
    .b(al_222a5f4d[33]),
    .c(al_222a5f4d[34]),
    .d(al_632b75dc[29]),
    .o(al_855effe8));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fea31acc (
    .a(al_855effe8),
    .b(al_4a463b38[27]),
    .c(al_632b75dc[24]),
    .o(al_e343d659[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2cab66c3 (
    .a(al_855effe8),
    .b(al_4a463b38[28]),
    .c(al_632b75dc[25]),
    .o(al_e343d659[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f4f4898a (
    .a(al_855effe8),
    .b(al_4a463b38[29]),
    .c(al_632b75dc[26]),
    .o(al_e343d659[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a7e1c26 (
    .a(al_855effe8),
    .b(al_4a463b38[30]),
    .c(al_632b75dc[27]),
    .o(al_e343d659[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b425bcf (
    .a(al_855effe8),
    .b(al_4a463b38[31]),
    .c(al_632b75dc[28]),
    .o(al_e343d659[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c864cb33 (
    .a(al_855effe8),
    .b(al_4a463b38[3]),
    .c(al_632b75dc[0]),
    .o(al_e343d659[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_607a2fe6 (
    .a(al_855effe8),
    .b(al_4a463b38[4]),
    .c(al_632b75dc[1]),
    .o(al_e343d659[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5b828d9e (
    .a(al_855effe8),
    .b(al_4a463b38[5]),
    .c(al_632b75dc[2]),
    .o(al_e343d659[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8f177908 (
    .a(al_855effe8),
    .b(al_4a463b38[6]),
    .c(al_632b75dc[3]),
    .o(al_e343d659[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a63b076 (
    .a(al_855effe8),
    .b(al_4a463b38[7]),
    .c(al_632b75dc[4]),
    .o(al_e343d659[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34cca471 (
    .a(al_855effe8),
    .b(al_4a463b38[8]),
    .c(al_632b75dc[5]),
    .o(al_e343d659[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93d72a0b (
    .a(al_855effe8),
    .b(al_4a463b38[9]),
    .c(al_632b75dc[6]),
    .o(al_e343d659[9]));
  AL_DFF_X al_1916d299 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0e2aae4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5db428bb[0]));
  AL_DFF_X al_c7056efe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[8]));
  AL_DFF_X al_10971f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[9]));
  AL_DFF_X al_a27a137 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[10]));
  AL_DFF_X al_fbe71f65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[11]));
  AL_DFF_X al_dcbb13d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[12]));
  AL_DFF_X al_72f2d76c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[13]));
  AL_DFF_X al_dad113ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[14]));
  AL_DFF_X al_b1f0c289 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[15]));
  AL_DFF_X al_af1a7c1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[16]));
  AL_DFF_X al_a419c583 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[17]));
  AL_DFF_X al_79515273 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[18]));
  AL_DFF_X al_db375e98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[19]));
  AL_DFF_X al_bc047058 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[20]));
  AL_DFF_X al_1e6ab7c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[21]));
  AL_DFF_X al_8c967d54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[22]));
  AL_DFF_X al_e201a3f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[23]));
  AL_DFF_X al_8e8e5f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[24]));
  AL_DFF_X al_4604158b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[25]));
  AL_DFF_X al_cf331084 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[26]));
  AL_DFF_X al_fc1dd323 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[27]));
  AL_DFF_X al_c2407fab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[28]));
  AL_DFF_X al_fd3268b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[29]));
  AL_DFF_X al_3426bb42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[30]));
  AL_DFF_X al_ca5ae43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[31]));
  AL_DFF_X al_aeb26b40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[32]));
  AL_DFF_X al_33a6761d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[33]));
  AL_DFF_X al_b24d2e93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[2]));
  AL_DFF_X al_1503a984 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[3]));
  AL_DFF_X al_eae81508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[4]));
  AL_DFF_X al_69e5a399 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[5]));
  AL_DFF_X al_264722a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[6]));
  AL_DFF_X al_2ecc103b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[7]));
  AL_DFF_X al_53d551bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[8]));
  AL_DFF_X al_faf5bbad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[9]));
  AL_DFF_X al_de49d4d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[10]));
  AL_DFF_X al_8e74d99a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[11]));
  AL_DFF_X al_4d28515c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[12]));
  AL_DFF_X al_3c0a6785 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[13]));
  AL_DFF_X al_540cd374 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[14]));
  AL_DFF_X al_545a6106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[15]));
  AL_DFF_X al_69a839f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[16]));
  AL_DFF_X al_3304dcb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[17]));
  AL_DFF_X al_ce1e62d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[0]));
  AL_DFF_X al_60c65214 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[18]));
  AL_DFF_X al_34a4719c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[19]));
  AL_DFF_X al_f3940230 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[20]));
  AL_DFF_X al_7d35f262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[21]));
  AL_DFF_X al_4bb11620 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[22]));
  AL_DFF_X al_fbf6879e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[23]));
  AL_DFF_X al_ce7f39ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[24]));
  AL_DFF_X al_e73248ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[25]));
  AL_DFF_X al_eec17c59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[26]));
  AL_DFF_X al_d66aa284 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[27]));
  AL_DFF_X al_be6e473b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[1]));
  AL_DFF_X al_a63cdb8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[28]));
  AL_DFF_X al_5b1245a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[29]));
  AL_DFF_X al_b1ae11f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[30]));
  AL_DFF_X al_66132836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[31]));
  AL_DFF_X al_599f62a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[2]));
  AL_DFF_X al_deac03ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[3]));
  AL_DFF_X al_6559dc3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[4]));
  AL_DFF_X al_c51e943b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[5]));
  AL_DFF_X al_4a87e4b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[6]));
  AL_DFF_X al_32ef0ceb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[7]));
  AL_DFF_X al_eccc4423 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[8]));
  AL_DFF_X al_fc736ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[9]));
  AL_DFF_X al_2992ad92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[10]));
  AL_DFF_X al_65315284 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[11]));
  AL_DFF_X al_7951b749 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[12]));
  AL_DFF_X al_38a3e380 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[13]));
  AL_DFF_X al_a12f847 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[14]));
  AL_DFF_X al_cae5449c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[15]));
  AL_DFF_X al_8b33cb5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[16]));
  AL_DFF_X al_20723779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[17]));
  AL_DFF_X al_e73c54fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_855effe8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[0]));
  AL_DFF_X al_ca81af0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[18]));
  AL_DFF_X al_2bf778e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[19]));
  AL_DFF_X al_ee1d0fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[20]));
  AL_DFF_X al_7718ed16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[21]));
  AL_DFF_X al_b08b1771 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[22]));
  AL_DFF_X al_8c72c6e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[23]));
  AL_DFF_X al_b9072722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[24]));
  AL_DFF_X al_42e1dbaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[25]));
  AL_DFF_X al_21a232b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[26]));
  AL_DFF_X al_ee5b0e69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[27]));
  AL_DFF_X al_6db59327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[1]));
  AL_DFF_X al_aa6812b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[28]));
  AL_DFF_X al_8b3f1629 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[2]));
  AL_DFF_X al_ca0ece03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[3]));
  AL_DFF_X al_73d8b0d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[4]));
  AL_DFF_X al_73cee2b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[5]));
  AL_DFF_X al_f9400736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[6]));
  AL_DFF_X al_b3d5907 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_57399a9 (
    .a(1'b0),
    .o({al_966d3a1d,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ffb5771 (
    .a(al_32ba5b24[2]),
    .b(al_d1a07609[2]),
    .c(al_966d3a1d),
    .o({al_f4c9a2d4,al_10f8c714[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8711c39 (
    .a(al_32ba5b24[3]),
    .b(al_d1a07609[3]),
    .c(al_f4c9a2d4),
    .o({al_42dadf79,al_10f8c714[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_407df837 (
    .a(al_32ba5b24[4]),
    .b(al_d1a07609[4]),
    .c(al_42dadf79),
    .o({al_97bfe275,al_10f8c714[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13daa0bd (
    .a(al_32ba5b24[5]),
    .b(al_d1a07609[5]),
    .c(al_97bfe275),
    .o({al_8ef4e9d1,al_10f8c714[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bdb5f146 (
    .a(al_32ba5b24[6]),
    .b(al_d1a07609[6]),
    .c(al_8ef4e9d1),
    .o({al_1a4fdc2c,al_10f8c714[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7febb2a5 (
    .a(al_32ba5b24[7]),
    .b(al_d1a07609[7]),
    .c(al_1a4fdc2c),
    .o({al_99c43840,al_10f8c714[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8fcdff7d (
    .a(al_32ba5b24[8]),
    .b(al_d1a07609[8]),
    .c(al_99c43840),
    .o({al_98c65d85,al_10f8c714[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e899ce4 (
    .a(al_32ba5b24[9]),
    .b(al_d1a07609[9]),
    .c(al_98c65d85),
    .o({al_5b6cf04f,al_10f8c714[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c417cdf (
    .a(al_32ba5b24[10]),
    .b(al_d1a07609[10]),
    .c(al_5b6cf04f),
    .o({al_ae08306c,al_10f8c714[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8e020320 (
    .a(al_32ba5b24[11]),
    .b(al_d1a07609[11]),
    .c(al_ae08306c),
    .o({al_7f4546cf,al_10f8c714[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_62a2dafd (
    .a(al_32ba5b24[12]),
    .b(al_d1a07609[12]),
    .c(al_7f4546cf),
    .o({al_f23b4ac3,al_10f8c714[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9064caf9 (
    .a(al_32ba5b24[13]),
    .b(al_d1a07609[13]),
    .c(al_f23b4ac3),
    .o({al_ac9e4212,al_10f8c714[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_121b91a (
    .a(al_32ba5b24[14]),
    .b(al_d1a07609[14]),
    .c(al_ac9e4212),
    .o({al_78275fb6,al_10f8c714[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_93d24064 (
    .a(al_32ba5b24[15]),
    .b(al_d1a07609[15]),
    .c(al_78275fb6),
    .o({al_9a080fbf,al_10f8c714[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a8fbd71 (
    .a(al_32ba5b24[16]),
    .b(al_d1a07609[16]),
    .c(al_9a080fbf),
    .o({al_8a23505f,al_10f8c714[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f9982892 (
    .a(al_32ba5b24[17]),
    .b(al_d1a07609[17]),
    .c(al_8a23505f),
    .o({al_5f9068e6,al_10f8c714[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d78395 (
    .a(al_32ba5b24[18]),
    .b(al_d1a07609[18]),
    .c(al_5f9068e6),
    .o({al_a46f14d2,al_10f8c714[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dea27c86 (
    .a(al_32ba5b24[19]),
    .b(al_d1a07609[19]),
    .c(al_a46f14d2),
    .o({al_342b0ff9,al_10f8c714[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6fb58240 (
    .a(al_32ba5b24[20]),
    .b(al_d1a07609[20]),
    .c(al_342b0ff9),
    .o({al_e782992a,al_10f8c714[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84ba533c (
    .a(al_32ba5b24[21]),
    .b(al_d1a07609[21]),
    .c(al_e782992a),
    .o({al_5d589bca,al_10f8c714[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_11980c48 (
    .a(al_32ba5b24[22]),
    .b(al_d1a07609[22]),
    .c(al_5d589bca),
    .o({al_33f64520,al_10f8c714[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_100fe815 (
    .a(al_32ba5b24[23]),
    .b(al_d1a07609[23]),
    .c(al_33f64520),
    .o({al_e9c34253,al_10f8c714[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98d84602 (
    .a(al_32ba5b24[24]),
    .b(al_d1a07609[24]),
    .c(al_e9c34253),
    .o({al_d36ef0a6,al_10f8c714[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d82862c5 (
    .a(al_32ba5b24[25]),
    .b(al_d1a07609[25]),
    .c(al_d36ef0a6),
    .o({al_dd36b780,al_10f8c714[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7cbb4871 (
    .a(al_32ba5b24[26]),
    .b(al_d1a07609[26]),
    .c(al_dd36b780),
    .o({al_232ecfaf,al_10f8c714[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14f52b9a (
    .a(al_32ba5b24[27]),
    .b(al_d1a07609[27]),
    .c(al_232ecfaf),
    .o({al_f2fd9563,al_10f8c714[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b27244d (
    .a(al_32ba5b24[28]),
    .b(al_d1a07609[28]),
    .c(al_f2fd9563),
    .o({al_4c3e9ef3,al_10f8c714[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72937fea (
    .a(al_32ba5b24[29]),
    .b(al_d1a07609[29]),
    .c(al_4c3e9ef3),
    .o({al_6c944eaa,al_10f8c714[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7739c750 (
    .a(al_32ba5b24[30]),
    .b(al_d1a07609[30]),
    .c(al_6c944eaa),
    .o({al_8f677fc9,al_10f8c714[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9f0f19ad (
    .a(al_32ba5b24[31]),
    .b(al_d1a07609[31]),
    .c(al_8f677fc9),
    .o({al_5fcd8d3b,al_10f8c714[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_69f15862 (
    .c(al_5fcd8d3b),
    .o({open_n119,al_10f8c714[30]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_887708b1 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[10]),
    .c(al_10f8c714[8]),
    .o(al_14165a56[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_231f946 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[11]),
    .c(al_10f8c714[9]),
    .o(al_14165a56[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_89e9a643 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[12]),
    .c(al_10f8c714[10]),
    .o(al_14165a56[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d278bb24 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[13]),
    .c(al_10f8c714[11]),
    .o(al_14165a56[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_25c712f3 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[14]),
    .c(al_10f8c714[12]),
    .o(al_14165a56[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bc80b81e (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[15]),
    .c(al_10f8c714[13]),
    .o(al_14165a56[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b1009d6e (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[16]),
    .c(al_10f8c714[14]),
    .o(al_14165a56[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7fca3ef1 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[17]),
    .c(al_10f8c714[15]),
    .o(al_14165a56[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_239f1f05 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[18]),
    .c(al_10f8c714[16]),
    .o(al_14165a56[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c07aa2d5 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[19]),
    .c(al_10f8c714[17]),
    .o(al_14165a56[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f445c83 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[20]),
    .c(al_10f8c714[18]),
    .o(al_14165a56[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_caf5d5cc (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[21]),
    .c(al_10f8c714[19]),
    .o(al_14165a56[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1769f616 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[22]),
    .c(al_10f8c714[20]),
    .o(al_14165a56[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c92af4d (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[23]),
    .c(al_10f8c714[21]),
    .o(al_14165a56[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8a1fbdd (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[24]),
    .c(al_10f8c714[22]),
    .o(al_14165a56[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e8a834a0 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[25]),
    .c(al_10f8c714[23]),
    .o(al_14165a56[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_50cbb86b (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[26]),
    .c(al_10f8c714[24]),
    .o(al_14165a56[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f80656e (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[27]),
    .c(al_10f8c714[25]),
    .o(al_14165a56[27]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_e98bab02 (
    .a(al_d1a07609[32]),
    .b(al_d1a07609[33]),
    .c(al_10f8c714[30]),
    .o(al_5fd9abe8));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c6e86ff4 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[28]),
    .c(al_10f8c714[26]),
    .o(al_14165a56[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6080847d (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[29]),
    .c(al_10f8c714[27]),
    .o(al_14165a56[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_76cb45ff (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[2]),
    .c(al_10f8c714[0]),
    .o(al_14165a56[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4209a834 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[30]),
    .c(al_10f8c714[28]),
    .o(al_14165a56[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ddfa8cc3 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[31]),
    .c(al_10f8c714[29]),
    .o(al_14165a56[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e14347b9 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[3]),
    .c(al_10f8c714[1]),
    .o(al_14165a56[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ae67b63c (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[4]),
    .c(al_10f8c714[2]),
    .o(al_14165a56[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e80f9534 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[5]),
    .c(al_10f8c714[3]),
    .o(al_14165a56[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_17697983 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[6]),
    .c(al_10f8c714[4]),
    .o(al_14165a56[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_79045d50 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[7]),
    .c(al_10f8c714[5]),
    .o(al_14165a56[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_89a85ed6 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[8]),
    .c(al_10f8c714[6]),
    .o(al_14165a56[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7b833d4 (
    .a(al_5fd9abe8),
    .b(al_32ba5b24[9]),
    .c(al_10f8c714[7]),
    .o(al_14165a56[9]));
  AL_DFF_X al_7bac587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5db428bb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d805738[0]));
  AL_DFF_X al_8e895fb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[8]));
  AL_DFF_X al_6a1ed9ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[9]));
  AL_DFF_X al_a0ef1afb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[10]));
  AL_DFF_X al_cfe80524 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[11]));
  AL_DFF_X al_d63233bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[12]));
  AL_DFF_X al_83ea5181 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[13]));
  AL_DFF_X al_27910570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[14]));
  AL_DFF_X al_2f64d09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[15]));
  AL_DFF_X al_7782e3ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[16]));
  AL_DFF_X al_867a77db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[17]));
  AL_DFF_X al_b1a8552d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[18]));
  AL_DFF_X al_e509198b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[19]));
  AL_DFF_X al_ba8a655b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[20]));
  AL_DFF_X al_b0469ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[21]));
  AL_DFF_X al_e1cbbe41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[22]));
  AL_DFF_X al_3cda224a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[23]));
  AL_DFF_X al_30e89bcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[24]));
  AL_DFF_X al_72650096 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[25]));
  AL_DFF_X al_a7eb2eb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[26]));
  AL_DFF_X al_2004ff65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[27]));
  AL_DFF_X al_85ad7f97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[1]));
  AL_DFF_X al_18eb0ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[28]));
  AL_DFF_X al_25f3ec55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[29]));
  AL_DFF_X al_8c93f665 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[30]));
  AL_DFF_X al_d8f72f3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[31]));
  AL_DFF_X al_a2f3d7c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[32]));
  AL_DFF_X al_edac6efc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[2]));
  AL_DFF_X al_3aecd42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[3]));
  AL_DFF_X al_db21e8f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[4]));
  AL_DFF_X al_3a70a7ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[5]));
  AL_DFF_X al_928fc59a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[6]));
  AL_DFF_X al_7dcf84e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[7]));
  AL_DFF_X al_b35e3a94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[8]));
  AL_DFF_X al_762b7c06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[9]));
  AL_DFF_X al_99bffd28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[10]));
  AL_DFF_X al_90c8f5b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[11]));
  AL_DFF_X al_52eb3cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[12]));
  AL_DFF_X al_ac7ceb7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[13]));
  AL_DFF_X al_462d4ddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[14]));
  AL_DFF_X al_97a374f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[15]));
  AL_DFF_X al_c274eda6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[16]));
  AL_DFF_X al_fda9f5ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[17]));
  AL_DFF_X al_9e50d7cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[0]));
  AL_DFF_X al_9f68cc2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[18]));
  AL_DFF_X al_96c2fd9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[19]));
  AL_DFF_X al_a6babeb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[20]));
  AL_DFF_X al_14b01f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[21]));
  AL_DFF_X al_d778b855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[22]));
  AL_DFF_X al_7cc985ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[23]));
  AL_DFF_X al_7588bd8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[24]));
  AL_DFF_X al_f78868cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[25]));
  AL_DFF_X al_b0d0b537 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[26]));
  AL_DFF_X al_9832e889 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[27]));
  AL_DFF_X al_84fc67fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[1]));
  AL_DFF_X al_96976b89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[28]));
  AL_DFF_X al_f747906c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[29]));
  AL_DFF_X al_6347949c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[30]));
  AL_DFF_X al_70133822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[31]));
  AL_DFF_X al_81d4f594 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[2]));
  AL_DFF_X al_ef9a2c60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[3]));
  AL_DFF_X al_fed989ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[4]));
  AL_DFF_X al_b62c4cbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[5]));
  AL_DFF_X al_f741e71f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[6]));
  AL_DFF_X al_20cbe7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[7]));
  AL_DFF_X al_fc4b7e5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[8]));
  AL_DFF_X al_fd95e1d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[9]));
  AL_DFF_X al_2119bac6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[10]));
  AL_DFF_X al_ada85597 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[11]));
  AL_DFF_X al_6090af49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[12]));
  AL_DFF_X al_8f9f67d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[13]));
  AL_DFF_X al_f1bd1f59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[14]));
  AL_DFF_X al_b20b8242 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[15]));
  AL_DFF_X al_6e379f82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[16]));
  AL_DFF_X al_633f4270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[17]));
  AL_DFF_X al_66cdbd2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd9abe8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[0]));
  AL_DFF_X al_e448e50f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[18]));
  AL_DFF_X al_a5d9eec9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[19]));
  AL_DFF_X al_4d34e407 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[20]));
  AL_DFF_X al_7362068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[21]));
  AL_DFF_X al_ab3ba732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[22]));
  AL_DFF_X al_6f247955 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[23]));
  AL_DFF_X al_535f6d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[24]));
  AL_DFF_X al_8ec6b0b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[25]));
  AL_DFF_X al_9d6dc5ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[26]));
  AL_DFF_X al_eca54707 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[27]));
  AL_DFF_X al_6f0d0865 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[1]));
  AL_DFF_X al_88f060a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[28]));
  AL_DFF_X al_d0cc55db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[29]));
  AL_DFF_X al_d2012e87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[2]));
  AL_DFF_X al_c7357867 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[3]));
  AL_DFF_X al_1097e039 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[4]));
  AL_DFF_X al_b379612e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[5]));
  AL_DFF_X al_222a3732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[6]));
  AL_DFF_X al_1ee503a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_40b32c7b (
    .a(al_78d777d2),
    .b(al_853654c1),
    .c(al_5173861b),
    .o(al_7a77d617));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2aa166f (
    .a(al_6a637a32[48]),
    .b(al_6a637a32[49]),
    .c(al_6a637a32[50]),
    .d(al_6a637a32[51]),
    .e(al_6a637a32[52]),
    .f(al_6a637a32[53]),
    .o(al_56a083ea));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_9491b318 (
    .a(al_6a637a32[38]),
    .b(al_6a637a32[39]),
    .c(al_6a637a32[40]),
    .d(al_6a637a32[41]),
    .o(al_249d4728));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_97c28cec (
    .a(al_6769a627),
    .b(al_249d4728),
    .c(al_6a637a32[36]),
    .d(al_6a637a32[37]),
    .e(al_6a637a32[42]),
    .f(al_6a637a32[43]),
    .o(al_853654c1));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    .INIT(16'hf731))
    al_69beed7 (
    .a(al_6a637a32[29]),
    .b(al_6a637a32[30]),
    .c(al_3d0cfeb4[29]),
    .d(al_3d0cfeb4[30]),
    .o(al_6c21e4f));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*B*C)"),
    .INIT(8'h4d))
    al_880216bf (
    .a(al_6c21e4f),
    .b(al_6a637a32[31]),
    .c(al_3d0cfeb4[31]),
    .o(al_5173861b));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~C*B*A))"),
    .INIT(32'hf7ff0800))
    al_cc2a2a01 (
    .a(al_78d777d2),
    .b(al_853654c1),
    .c(al_5173861b),
    .d(al_6a637a32[29]),
    .e(al_3d0cfeb4[29]),
    .o(al_a9b28455[29]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_dbf5ee3c (
    .a(al_6a637a32[32]),
    .b(al_6a637a32[33]),
    .c(al_6a637a32[34]),
    .d(al_6a637a32[35]),
    .e(al_6a637a32[60]),
    .o(al_7028725));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3a23f591 (
    .a(al_6a637a32[56]),
    .b(al_6a637a32[57]),
    .c(al_6a637a32[58]),
    .d(al_6a637a32[59]),
    .o(al_aa188274));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_6bf9536d (
    .a(al_56a083ea),
    .b(al_7028725),
    .c(al_aa188274),
    .d(al_6a637a32[54]),
    .e(al_6a637a32[55]),
    .o(al_78d777d2));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7737ebbf (
    .a(al_6a637a32[44]),
    .b(al_6a637a32[45]),
    .c(al_6a637a32[46]),
    .d(al_6a637a32[47]),
    .o(al_6769a627));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*A))"),
    .INIT(8'hc6))
    al_3259f828 (
    .a(al_6a637a32[29]),
    .b(al_6a637a32[30]),
    .c(al_3d0cfeb4[29]),
    .o(al_1a0f9e95));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~C*B*A))"),
    .INIT(32'hf7ff0800))
    al_e492e415 (
    .a(al_78d777d2),
    .b(al_853654c1),
    .c(al_5173861b),
    .d(al_1a0f9e95),
    .e(al_3d0cfeb4[30]),
    .o(al_a9b28455[30]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(B*A*~(D@C)))"),
    .INIT(32'h7ff70000))
    al_40580873 (
    .a(al_78d777d2),
    .b(al_853654c1),
    .c(al_6c21e4f),
    .d(al_6a637a32[31]),
    .e(al_3d0cfeb4[31]),
    .o(al_a9b28455[31]));
  AL_DFF_X al_a3f6140e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_67f5b0b3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44882eca[0]));
  AL_DFF_X al_26872ba6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[28]));
  AL_DFF_X al_769c4989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[29]));
  AL_DFF_X al_ece0d1fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[30]));
  AL_DFF_X al_974aa297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[31]));
  AL_DFF_X al_3408a219 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[32]));
  AL_DFF_X al_d72283d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[33]));
  AL_DFF_X al_cecd4b01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[34]));
  AL_DFF_X al_b308f973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[35]));
  AL_DFF_X al_7c2ca730 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[36]));
  AL_DFF_X al_cfa06733 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[37]));
  AL_DFF_X al_238e5e1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[38]));
  AL_DFF_X al_c1bd4df7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[39]));
  AL_DFF_X al_3e038591 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[40]));
  AL_DFF_X al_13c9827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[41]));
  AL_DFF_X al_18e97e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[42]));
  AL_DFF_X al_ebd49d44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[43]));
  AL_DFF_X al_5fae692b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[44]));
  AL_DFF_X al_e63afd48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[45]));
  AL_DFF_X al_52898fd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[46]));
  AL_DFF_X al_a549dadf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[47]));
  AL_DFF_X al_5093188 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[48]));
  AL_DFF_X al_d633e346 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[49]));
  AL_DFF_X al_c2767705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[50]));
  AL_DFF_X al_e2b6799d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[51]));
  AL_DFF_X al_7bd5a7d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[52]));
  AL_DFF_X al_5bf9b570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[53]));
  AL_DFF_X al_9c5bdeff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[54]));
  AL_DFF_X al_15a6529e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[55]));
  AL_DFF_X al_ae273c16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[56]));
  AL_DFF_X al_d22ae3b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[57]));
  AL_DFF_X al_a76a94ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[58]));
  AL_DFF_X al_7ddb78b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[59]));
  AL_DFF_X al_eb6810df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[8]));
  AL_DFF_X al_660f57cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[9]));
  AL_DFF_X al_a14688f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[10]));
  AL_DFF_X al_16384734 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[11]));
  AL_DFF_X al_a81439c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[12]));
  AL_DFF_X al_eb8e93aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[13]));
  AL_DFF_X al_35eb088a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[14]));
  AL_DFF_X al_59059b2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[15]));
  AL_DFF_X al_6edec2f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[16]));
  AL_DFF_X al_e014fa3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[17]));
  AL_DFF_X al_19caaf92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[0]));
  AL_DFF_X al_685b63ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[18]));
  AL_DFF_X al_75d4ebb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[19]));
  AL_DFF_X al_8ece4b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[20]));
  AL_DFF_X al_af8ce59b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[21]));
  AL_DFF_X al_95f2b96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[22]));
  AL_DFF_X al_ef02eff6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[23]));
  AL_DFF_X al_db293ec9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[24]));
  AL_DFF_X al_8ef5c889 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[25]));
  AL_DFF_X al_1581088a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[26]));
  AL_DFF_X al_b18d6448 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[27]));
  AL_DFF_X al_4f1e9f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[1]));
  AL_DFF_X al_69df85fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[28]));
  AL_DFF_X al_f7005208 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[29]));
  AL_DFF_X al_da3742de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[30]));
  AL_DFF_X al_da94f051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[31]));
  AL_DFF_X al_f8d428bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[2]));
  AL_DFF_X al_68091650 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[3]));
  AL_DFF_X al_e2810320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[4]));
  AL_DFF_X al_7c1769ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[5]));
  AL_DFF_X al_6c250488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[6]));
  AL_DFF_X al_c179f202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[7]));
  AL_DFF_X al_ee02adcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a77d617),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[0]));
  AL_DFF_X al_143a9a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b54c1014[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[1]));
  AL_DFF_X al_f44364e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b54c1014[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[2]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_152cce9e (
    .a(1'b0),
    .o({al_4f5a23d4,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_739dba21 (
    .a(al_690b21a4[1]),
    .b(al_627988c3[1]),
    .c(al_4f5a23d4),
    .o({al_3eebd40f,al_7c1783ce[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d3a8c26d (
    .a(al_690b21a4[2]),
    .b(al_627988c3[2]),
    .c(al_3eebd40f),
    .o({al_8e4361ca,al_7c1783ce[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92eeb4c5 (
    .a(al_690b21a4[3]),
    .b(al_627988c3[3]),
    .c(al_8e4361ca),
    .o({al_912de09d,al_7c1783ce[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14e762d3 (
    .a(al_690b21a4[4]),
    .b(al_627988c3[4]),
    .c(al_912de09d),
    .o({al_85cca751,al_7c1783ce[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9a8b9d2 (
    .a(al_690b21a4[5]),
    .b(al_627988c3[5]),
    .c(al_85cca751),
    .o({al_ad8d6e84,al_7c1783ce[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_56cf2b39 (
    .a(al_690b21a4[6]),
    .b(al_627988c3[6]),
    .c(al_ad8d6e84),
    .o({al_5992e66f,al_7c1783ce[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a15876a7 (
    .a(al_690b21a4[7]),
    .b(al_627988c3[7]),
    .c(al_5992e66f),
    .o({al_53645fd3,al_7c1783ce[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f82256a (
    .a(al_690b21a4[8]),
    .b(al_627988c3[8]),
    .c(al_53645fd3),
    .o({al_5c00f664,al_7c1783ce[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e791ad44 (
    .a(al_690b21a4[9]),
    .b(al_627988c3[9]),
    .c(al_5c00f664),
    .o({al_a5fb5d66,al_7c1783ce[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_352d30a1 (
    .a(al_690b21a4[10]),
    .b(al_627988c3[10]),
    .c(al_a5fb5d66),
    .o({al_bfb57bee,al_7c1783ce[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d16d4f29 (
    .a(al_690b21a4[11]),
    .b(al_627988c3[11]),
    .c(al_bfb57bee),
    .o({al_2f85c10c,al_7c1783ce[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_29064497 (
    .a(al_690b21a4[12]),
    .b(al_627988c3[12]),
    .c(al_2f85c10c),
    .o({al_ce21f8f3,al_7c1783ce[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a5f7538c (
    .a(al_690b21a4[13]),
    .b(al_627988c3[13]),
    .c(al_ce21f8f3),
    .o({al_83736e7b,al_7c1783ce[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a741b0dd (
    .a(al_690b21a4[14]),
    .b(al_627988c3[14]),
    .c(al_83736e7b),
    .o({al_c3f591aa,al_7c1783ce[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8627535f (
    .a(al_690b21a4[15]),
    .b(al_627988c3[15]),
    .c(al_c3f591aa),
    .o({al_fbb0bdd6,al_7c1783ce[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_863928d8 (
    .a(al_690b21a4[16]),
    .b(al_627988c3[16]),
    .c(al_fbb0bdd6),
    .o({al_eb11562b,al_7c1783ce[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a2c376 (
    .a(al_690b21a4[17]),
    .b(al_627988c3[17]),
    .c(al_eb11562b),
    .o({al_15d2d0ed,al_7c1783ce[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36176996 (
    .a(al_690b21a4[18]),
    .b(al_627988c3[18]),
    .c(al_15d2d0ed),
    .o({al_a792d40a,al_7c1783ce[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cce2f41e (
    .a(al_690b21a4[19]),
    .b(al_627988c3[19]),
    .c(al_a792d40a),
    .o({al_92024dcf,al_7c1783ce[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9a4d29f2 (
    .a(al_690b21a4[20]),
    .b(al_627988c3[20]),
    .c(al_92024dcf),
    .o({al_60518bd5,al_7c1783ce[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d94cc882 (
    .a(al_690b21a4[21]),
    .b(al_627988c3[21]),
    .c(al_60518bd5),
    .o({al_a0662365,al_7c1783ce[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_22d84dc2 (
    .a(al_690b21a4[22]),
    .b(al_627988c3[22]),
    .c(al_a0662365),
    .o({al_d44591b2,al_7c1783ce[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_896fe8e9 (
    .a(al_690b21a4[23]),
    .b(al_627988c3[23]),
    .c(al_d44591b2),
    .o({al_1280dac2,al_7c1783ce[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfee239 (
    .a(al_690b21a4[24]),
    .b(al_627988c3[24]),
    .c(al_1280dac2),
    .o({al_655899d3,al_7c1783ce[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1a618971 (
    .a(al_690b21a4[25]),
    .b(al_627988c3[25]),
    .c(al_655899d3),
    .o({al_3a98aee3,al_7c1783ce[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8753718 (
    .a(al_690b21a4[26]),
    .b(al_627988c3[26]),
    .c(al_3a98aee3),
    .o({al_6269677,al_7c1783ce[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13dd7485 (
    .a(al_690b21a4[27]),
    .b(al_627988c3[27]),
    .c(al_6269677),
    .o({al_f6aa030f,al_7c1783ce[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_707dd93a (
    .a(al_690b21a4[28]),
    .b(al_627988c3[28]),
    .c(al_f6aa030f),
    .o({al_1e3baa15,al_7c1783ce[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a65264e5 (
    .a(al_690b21a4[29]),
    .b(al_627988c3[29]),
    .c(al_1e3baa15),
    .o({al_90c4774,al_7c1783ce[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a383a976 (
    .a(al_690b21a4[30]),
    .b(al_627988c3[30]),
    .c(al_90c4774),
    .o({al_2d7cd5be,al_7c1783ce[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8e9ecbb4 (
    .a(al_690b21a4[31]),
    .b(al_627988c3[31]),
    .c(al_2d7cd5be),
    .o({al_41002c4f,al_7c1783ce[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f9a9dfb6 (
    .c(al_41002c4f),
    .o({open_n125,al_7c1783ce[31]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_453f2889 (
    .a(al_b06c909),
    .b(al_690b21a4[10]),
    .c(al_7c1783ce[9]),
    .o(al_3ccb3a4f[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7e04688f (
    .a(al_b06c909),
    .b(al_690b21a4[11]),
    .c(al_7c1783ce[10]),
    .o(al_3ccb3a4f[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99d5a0ec (
    .a(al_b06c909),
    .b(al_690b21a4[12]),
    .c(al_7c1783ce[11]),
    .o(al_3ccb3a4f[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8091872d (
    .a(al_b06c909),
    .b(al_690b21a4[13]),
    .c(al_7c1783ce[12]),
    .o(al_3ccb3a4f[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3e3bd2b (
    .a(al_b06c909),
    .b(al_690b21a4[14]),
    .c(al_7c1783ce[13]),
    .o(al_3ccb3a4f[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b3b54b04 (
    .a(al_b06c909),
    .b(al_690b21a4[15]),
    .c(al_7c1783ce[14]),
    .o(al_3ccb3a4f[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c6d7974 (
    .a(al_b06c909),
    .b(al_690b21a4[16]),
    .c(al_7c1783ce[15]),
    .o(al_3ccb3a4f[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_971e1476 (
    .a(al_b06c909),
    .b(al_690b21a4[17]),
    .c(al_7c1783ce[16]),
    .o(al_3ccb3a4f[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_912b0dd0 (
    .a(al_b06c909),
    .b(al_690b21a4[18]),
    .c(al_7c1783ce[17]),
    .o(al_3ccb3a4f[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da7f19aa (
    .a(al_b06c909),
    .b(al_690b21a4[19]),
    .c(al_7c1783ce[18]),
    .o(al_3ccb3a4f[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93be6fc8 (
    .a(al_b06c909),
    .b(al_690b21a4[1]),
    .c(al_7c1783ce[0]),
    .o(al_3ccb3a4f[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_329f04d4 (
    .a(al_b06c909),
    .b(al_690b21a4[20]),
    .c(al_7c1783ce[19]),
    .o(al_3ccb3a4f[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_38fb5244 (
    .a(al_b06c909),
    .b(al_690b21a4[21]),
    .c(al_7c1783ce[20]),
    .o(al_3ccb3a4f[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b77668a5 (
    .a(al_b06c909),
    .b(al_690b21a4[22]),
    .c(al_7c1783ce[21]),
    .o(al_3ccb3a4f[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b0a229ca (
    .a(al_b06c909),
    .b(al_690b21a4[23]),
    .c(al_7c1783ce[22]),
    .o(al_3ccb3a4f[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f62d7f63 (
    .a(al_b06c909),
    .b(al_690b21a4[24]),
    .c(al_7c1783ce[23]),
    .o(al_3ccb3a4f[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7583c301 (
    .a(al_b06c909),
    .b(al_690b21a4[25]),
    .c(al_7c1783ce[24]),
    .o(al_3ccb3a4f[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_505a1d48 (
    .a(al_b06c909),
    .b(al_690b21a4[26]),
    .c(al_7c1783ce[25]),
    .o(al_3ccb3a4f[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bd67a4d5 (
    .a(al_b06c909),
    .b(al_690b21a4[27]),
    .c(al_7c1783ce[26]),
    .o(al_3ccb3a4f[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9d2c0b95 (
    .a(al_b06c909),
    .b(al_690b21a4[28]),
    .c(al_7c1783ce[27]),
    .o(al_3ccb3a4f[28]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_667996f6 (
    .a(al_627988c3[32]),
    .b(al_7c1783ce[31]),
    .o(al_b06c909));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8a73c4a5 (
    .a(al_b06c909),
    .b(al_690b21a4[29]),
    .c(al_7c1783ce[28]),
    .o(al_3ccb3a4f[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_830aef5f (
    .a(al_b06c909),
    .b(al_690b21a4[2]),
    .c(al_7c1783ce[1]),
    .o(al_3ccb3a4f[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9e4c789e (
    .a(al_b06c909),
    .b(al_690b21a4[30]),
    .c(al_7c1783ce[29]),
    .o(al_3ccb3a4f[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f4400b70 (
    .a(al_b06c909),
    .b(al_690b21a4[31]),
    .c(al_7c1783ce[30]),
    .o(al_3ccb3a4f[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f031819 (
    .a(al_b06c909),
    .b(al_690b21a4[3]),
    .c(al_7c1783ce[2]),
    .o(al_3ccb3a4f[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2a144a62 (
    .a(al_b06c909),
    .b(al_690b21a4[4]),
    .c(al_7c1783ce[3]),
    .o(al_3ccb3a4f[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a2e772be (
    .a(al_b06c909),
    .b(al_690b21a4[5]),
    .c(al_7c1783ce[4]),
    .o(al_3ccb3a4f[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_240b55a (
    .a(al_b06c909),
    .b(al_690b21a4[6]),
    .c(al_7c1783ce[5]),
    .o(al_3ccb3a4f[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ebd16b62 (
    .a(al_b06c909),
    .b(al_690b21a4[7]),
    .c(al_7c1783ce[6]),
    .o(al_3ccb3a4f[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9ab9aad9 (
    .a(al_b06c909),
    .b(al_690b21a4[8]),
    .c(al_7c1783ce[7]),
    .o(al_3ccb3a4f[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_579c78f1 (
    .a(al_b06c909),
    .b(al_690b21a4[9]),
    .c(al_7c1783ce[8]),
    .o(al_3ccb3a4f[9]));
  AL_DFF_X al_75205bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d805738[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74993dd2[0]));
  AL_DFF_X al_48129714 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[8]));
  AL_DFF_X al_3b315749 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[9]));
  AL_DFF_X al_5a83e029 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[10]));
  AL_DFF_X al_94ea4b89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[11]));
  AL_DFF_X al_3d3f59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[12]));
  AL_DFF_X al_4f82ddfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[13]));
  AL_DFF_X al_896a5c0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[14]));
  AL_DFF_X al_f77ddae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[15]));
  AL_DFF_X al_43edbfdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[16]));
  AL_DFF_X al_44adae8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[17]));
  AL_DFF_X al_5824b41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[0]));
  AL_DFF_X al_ba19e94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[18]));
  AL_DFF_X al_7059f920 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[19]));
  AL_DFF_X al_50e27670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[20]));
  AL_DFF_X al_279a4eaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[21]));
  AL_DFF_X al_b799be1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[22]));
  AL_DFF_X al_e11cbbec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[23]));
  AL_DFF_X al_2196b19b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[24]));
  AL_DFF_X al_7d10f985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[25]));
  AL_DFF_X al_cfdf44d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[26]));
  AL_DFF_X al_53b6cb78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[27]));
  AL_DFF_X al_5609839f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[1]));
  AL_DFF_X al_b29221f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[28]));
  AL_DFF_X al_cb296a2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[29]));
  AL_DFF_X al_759629b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[30]));
  AL_DFF_X al_92ff6e83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[31]));
  AL_DFF_X al_f3bf9e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[2]));
  AL_DFF_X al_80e9948c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[3]));
  AL_DFF_X al_1bca6ab1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[4]));
  AL_DFF_X al_d0b9ab9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[5]));
  AL_DFF_X al_d1ade42d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[6]));
  AL_DFF_X al_3d03f0ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[7]));
  AL_DFF_X al_90d96ad0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[8]));
  AL_DFF_X al_59877554 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[9]));
  AL_DFF_X al_1611287d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[10]));
  AL_DFF_X al_f09e7e10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[11]));
  AL_DFF_X al_67d7bbfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[12]));
  AL_DFF_X al_6103e1c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[13]));
  AL_DFF_X al_c6fb8ffe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[14]));
  AL_DFF_X al_c8b11b8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[15]));
  AL_DFF_X al_60a53f9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[16]));
  AL_DFF_X al_e9914b84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[17]));
  AL_DFF_X al_b861af81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[0]));
  AL_DFF_X al_ffba9671 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[18]));
  AL_DFF_X al_95a79d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[19]));
  AL_DFF_X al_96b7aee8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[20]));
  AL_DFF_X al_505cd9d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[21]));
  AL_DFF_X al_a526ff9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[22]));
  AL_DFF_X al_1b758bed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[23]));
  AL_DFF_X al_3c4efe7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[24]));
  AL_DFF_X al_8902aed2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[25]));
  AL_DFF_X al_ba16ebb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[26]));
  AL_DFF_X al_4cf25401 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[27]));
  AL_DFF_X al_2c70f2e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[1]));
  AL_DFF_X al_16cd9134 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[28]));
  AL_DFF_X al_7dcddf30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[29]));
  AL_DFF_X al_9cb18fa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[30]));
  AL_DFF_X al_cd11e96f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[31]));
  AL_DFF_X al_5f71c232 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[2]));
  AL_DFF_X al_8a93d8bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[3]));
  AL_DFF_X al_2188eeb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[4]));
  AL_DFF_X al_3a473d66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[5]));
  AL_DFF_X al_4b52d994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[6]));
  AL_DFF_X al_25357512 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[7]));
  AL_DFF_X al_1337124d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[8]));
  AL_DFF_X al_324af66d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[9]));
  AL_DFF_X al_7524f1ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[10]));
  AL_DFF_X al_49cd264f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[11]));
  AL_DFF_X al_c6809b32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[12]));
  AL_DFF_X al_7b625971 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[13]));
  AL_DFF_X al_d8d56dd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[14]));
  AL_DFF_X al_d34378e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[15]));
  AL_DFF_X al_bd8d62e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[16]));
  AL_DFF_X al_6779f42c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[17]));
  AL_DFF_X al_4ed37a41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b06c909),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[0]));
  AL_DFF_X al_1c3ac839 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[18]));
  AL_DFF_X al_47c037f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[19]));
  AL_DFF_X al_b046f0f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[20]));
  AL_DFF_X al_90c98704 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[21]));
  AL_DFF_X al_791620db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[22]));
  AL_DFF_X al_22255e87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[23]));
  AL_DFF_X al_3f5fef52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[24]));
  AL_DFF_X al_fe4edd30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[25]));
  AL_DFF_X al_df52abc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[26]));
  AL_DFF_X al_afb243f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[27]));
  AL_DFF_X al_46930f39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[1]));
  AL_DFF_X al_a9e6309a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[28]));
  AL_DFF_X al_fe161876 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[29]));
  AL_DFF_X al_6d3bedfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[30]));
  AL_DFF_X al_39ca96a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[2]));
  AL_DFF_X al_c648a3fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[3]));
  AL_DFF_X al_4a4b2451 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[4]));
  AL_DFF_X al_420bcee8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[5]));
  AL_DFF_X al_42462a9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[6]));
  AL_DFF_X al_b3852f46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_67b37726 (
    .a(al_57dc9b0c[0]),
    .b(al_df3b43b5[0]),
    .c(al_42f85898),
    .o(al_eb7d14b9[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4819cb52 (
    .a(al_57dc9b0c[10]),
    .b(al_df3b43b5[10]),
    .c(al_42f85898),
    .o(al_eb7d14b9[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dacb2900 (
    .a(al_57dc9b0c[11]),
    .b(al_df3b43b5[11]),
    .c(al_42f85898),
    .o(al_eb7d14b9[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8d4289d4 (
    .a(al_57dc9b0c[12]),
    .b(al_df3b43b5[12]),
    .c(al_42f85898),
    .o(al_eb7d14b9[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_435858ab (
    .a(al_57dc9b0c[13]),
    .b(al_df3b43b5[13]),
    .c(al_42f85898),
    .o(al_eb7d14b9[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bcbc9967 (
    .a(al_57dc9b0c[14]),
    .b(al_df3b43b5[14]),
    .c(al_42f85898),
    .o(al_eb7d14b9[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4145afa9 (
    .a(al_57dc9b0c[15]),
    .b(al_df3b43b5[15]),
    .c(al_42f85898),
    .o(al_eb7d14b9[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_48654d0a (
    .a(al_57dc9b0c[16]),
    .b(al_df3b43b5[16]),
    .c(al_42f85898),
    .o(al_eb7d14b9[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_42074f6b (
    .a(al_57dc9b0c[17]),
    .b(al_df3b43b5[17]),
    .c(al_42f85898),
    .o(al_eb7d14b9[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9aaf0dc1 (
    .a(al_57dc9b0c[18]),
    .b(al_df3b43b5[18]),
    .c(al_42f85898),
    .o(al_eb7d14b9[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8e71634d (
    .a(al_57dc9b0c[19]),
    .b(al_df3b43b5[19]),
    .c(al_42f85898),
    .o(al_eb7d14b9[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ba753ff5 (
    .a(al_57dc9b0c[1]),
    .b(al_df3b43b5[1]),
    .c(al_42f85898),
    .o(al_eb7d14b9[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6b7d1d91 (
    .a(al_57dc9b0c[20]),
    .b(al_df3b43b5[20]),
    .c(al_42f85898),
    .o(al_eb7d14b9[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c4ca852d (
    .a(al_57dc9b0c[21]),
    .b(al_df3b43b5[21]),
    .c(al_42f85898),
    .o(al_eb7d14b9[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4fbbad5a (
    .a(al_57dc9b0c[22]),
    .b(al_df3b43b5[22]),
    .c(al_42f85898),
    .o(al_eb7d14b9[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9439a588 (
    .a(al_57dc9b0c[23]),
    .b(al_df3b43b5[23]),
    .c(al_42f85898),
    .o(al_eb7d14b9[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_13239049 (
    .a(al_57dc9b0c[24]),
    .b(al_df3b43b5[24]),
    .c(al_42f85898),
    .o(al_eb7d14b9[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1c4c4b16 (
    .a(al_57dc9b0c[25]),
    .b(al_df3b43b5[25]),
    .c(al_42f85898),
    .o(al_eb7d14b9[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_84a0d2fc (
    .a(al_57dc9b0c[26]),
    .b(al_df3b43b5[26]),
    .c(al_42f85898),
    .o(al_eb7d14b9[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f7fb8903 (
    .a(al_57dc9b0c[27]),
    .b(al_df3b43b5[27]),
    .c(al_42f85898),
    .o(al_eb7d14b9[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_50f77443 (
    .a(al_57dc9b0c[28]),
    .b(al_df3b43b5[28]),
    .c(al_42f85898),
    .o(al_eb7d14b9[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ae46e3e5 (
    .a(al_57dc9b0c[29]),
    .b(al_df3b43b5[29]),
    .c(al_42f85898),
    .o(al_eb7d14b9[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fdbb6a37 (
    .a(al_57dc9b0c[2]),
    .b(al_df3b43b5[2]),
    .c(al_42f85898),
    .o(al_eb7d14b9[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ef45ea44 (
    .a(al_57dc9b0c[30]),
    .b(al_df3b43b5[30]),
    .c(al_42f85898),
    .o(al_eb7d14b9[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_216990ac (
    .a(al_57dc9b0c[31]),
    .b(al_df3b43b5[31]),
    .c(al_42f85898),
    .o(al_eb7d14b9[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_32295743 (
    .a(al_57dc9b0c[3]),
    .b(al_df3b43b5[3]),
    .c(al_42f85898),
    .o(al_eb7d14b9[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bb0502c1 (
    .a(al_57dc9b0c[4]),
    .b(al_df3b43b5[4]),
    .c(al_42f85898),
    .o(al_eb7d14b9[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6494fa40 (
    .a(al_57dc9b0c[5]),
    .b(al_df3b43b5[5]),
    .c(al_42f85898),
    .o(al_eb7d14b9[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cc190f2 (
    .a(al_57dc9b0c[6]),
    .b(al_df3b43b5[6]),
    .c(al_42f85898),
    .o(al_eb7d14b9[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e96b37e5 (
    .a(al_57dc9b0c[7]),
    .b(al_df3b43b5[7]),
    .c(al_42f85898),
    .o(al_eb7d14b9[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_260b607 (
    .a(al_57dc9b0c[8]),
    .b(al_df3b43b5[8]),
    .c(al_42f85898),
    .o(al_eb7d14b9[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f700e96f (
    .a(al_57dc9b0c[9]),
    .b(al_df3b43b5[9]),
    .c(al_42f85898),
    .o(al_eb7d14b9[9]));
  AL_DFF_X al_2e30312b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_74993dd2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5d831a[0]));
  AL_DFF_X al_2a4a0d84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[8]));
  AL_DFF_X al_ae1e8234 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[9]));
  AL_DFF_X al_eb0a6c18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[10]));
  AL_DFF_X al_d534ae55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[11]));
  AL_DFF_X al_7b990670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[12]));
  AL_DFF_X al_b1d4edb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[13]));
  AL_DFF_X al_61cb542d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[14]));
  AL_DFF_X al_d32f63a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[15]));
  AL_DFF_X al_1763af21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[16]));
  AL_DFF_X al_6b34549c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[17]));
  AL_DFF_X al_495ff80a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[0]));
  AL_DFF_X al_f3b299d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[18]));
  AL_DFF_X al_4295b698 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[19]));
  AL_DFF_X al_9b76de7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[20]));
  AL_DFF_X al_78450ef5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[21]));
  AL_DFF_X al_baf52ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[22]));
  AL_DFF_X al_42c4f73e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[23]));
  AL_DFF_X al_3bafea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[24]));
  AL_DFF_X al_973d97bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[25]));
  AL_DFF_X al_bc0e5550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[26]));
  AL_DFF_X al_61574c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[27]));
  AL_DFF_X al_c52346c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[1]));
  AL_DFF_X al_32c72431 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[28]));
  AL_DFF_X al_8783309e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[29]));
  AL_DFF_X al_c8f3dd9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[30]));
  AL_DFF_X al_a5e32e5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[31]));
  AL_DFF_X al_91a4d34f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[2]));
  AL_DFF_X al_ccdefea2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[3]));
  AL_DFF_X al_98c5dfdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[4]));
  AL_DFF_X al_40be9bd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[5]));
  AL_DFF_X al_41a25361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[6]));
  AL_DFF_X al_f65bab88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3519ff8d[7]));
  AL_DFF_X al_87fe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[8]));
  AL_DFF_X al_b3e960f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[9]));
  AL_DFF_X al_cedb61cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[10]));
  AL_DFF_X al_5f76df44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[11]));
  AL_DFF_X al_48f2f248 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[12]));
  AL_DFF_X al_971215ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[13]));
  AL_DFF_X al_fdbd2634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[14]));
  AL_DFF_X al_ea945541 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[15]));
  AL_DFF_X al_eca04bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[16]));
  AL_DFF_X al_75ebed64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[17]));
  AL_DFF_X al_65e79d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_42f85898),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[0]));
  AL_DFF_X al_72bf32af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[18]));
  AL_DFF_X al_247a9700 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[19]));
  AL_DFF_X al_98dae0e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[20]));
  AL_DFF_X al_df792ae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[21]));
  AL_DFF_X al_e9ff1687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[22]));
  AL_DFF_X al_be0492f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[23]));
  AL_DFF_X al_db20275a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[24]));
  AL_DFF_X al_33e8c553 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[25]));
  AL_DFF_X al_11580f51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[26]));
  AL_DFF_X al_2a719ef8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[27]));
  AL_DFF_X al_8a90b4e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[1]));
  AL_DFF_X al_e84fd4b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[28]));
  AL_DFF_X al_932b5679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[29]));
  AL_DFF_X al_a46a42d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[30]));
  AL_DFF_X al_a09b993d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[31]));
  AL_DFF_X al_62bb3fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[2]));
  AL_DFF_X al_5b7730d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[3]));
  AL_DFF_X al_96feeadc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[4]));
  AL_DFF_X al_bc902b89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[5]));
  AL_DFF_X al_727474fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[6]));
  AL_DFF_X al_1da0e0da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_18157fe8[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_576030d (
    .a(al_57dc9b0c[7]),
    .b(al_a5e9c08d[7]),
    .c(al_d720b206),
    .o({al_b05ac301,al_df3b43b5[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e4029bb (
    .a(al_57dc9b0c[8]),
    .b(al_a5e9c08d[8]),
    .c(al_b05ac301),
    .o({al_67046fd1,al_df3b43b5[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3e25337c (
    .a(al_57dc9b0c[9]),
    .b(al_a5e9c08d[9]),
    .c(al_67046fd1),
    .o({al_108156ff,al_df3b43b5[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a51b0652 (
    .a(al_57dc9b0c[10]),
    .b(al_a5e9c08d[10]),
    .c(al_108156ff),
    .o({al_162e0df5,al_df3b43b5[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de850a4b (
    .a(al_57dc9b0c[11]),
    .b(al_a5e9c08d[11]),
    .c(al_162e0df5),
    .o({al_61845f15,al_df3b43b5[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5033cba0 (
    .a(al_57dc9b0c[12]),
    .b(al_a5e9c08d[12]),
    .c(al_61845f15),
    .o({al_17de8af8,al_df3b43b5[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a22791c6 (
    .a(al_57dc9b0c[13]),
    .b(al_a5e9c08d[13]),
    .c(al_17de8af8),
    .o({al_e9f8df12,al_df3b43b5[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6eca77c1 (
    .a(al_57dc9b0c[14]),
    .b(al_a5e9c08d[14]),
    .c(al_e9f8df12),
    .o({al_e7a7f7d2,al_df3b43b5[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7956b96 (
    .a(al_57dc9b0c[15]),
    .b(al_a5e9c08d[15]),
    .c(al_e7a7f7d2),
    .o({al_37282f35,al_df3b43b5[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_919343b8 (
    .a(al_57dc9b0c[16]),
    .b(al_a5e9c08d[16]),
    .c(al_37282f35),
    .o({al_e1b1cb21,al_df3b43b5[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_bbc3ffe2 (
    .a(1'b0),
    .o({al_bb31a1fd,open_n128}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_811618a0 (
    .a(al_57dc9b0c[17]),
    .b(al_a5e9c08d[17]),
    .c(al_e1b1cb21),
    .o({al_eb87db38,al_df3b43b5[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3aa7ad7c (
    .a(al_57dc9b0c[18]),
    .b(al_a5e9c08d[18]),
    .c(al_eb87db38),
    .o({al_8db59e87,al_df3b43b5[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c4714d5d (
    .a(al_57dc9b0c[19]),
    .b(al_a5e9c08d[19]),
    .c(al_8db59e87),
    .o({al_8fa4d3c,al_df3b43b5[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_77f62dca (
    .a(al_57dc9b0c[20]),
    .b(al_a5e9c08d[20]),
    .c(al_8fa4d3c),
    .o({al_eddac2b0,al_df3b43b5[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_490553ef (
    .a(al_57dc9b0c[21]),
    .b(al_a5e9c08d[21]),
    .c(al_eddac2b0),
    .o({al_a23f6f13,al_df3b43b5[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1cdf1331 (
    .a(al_57dc9b0c[22]),
    .b(al_a5e9c08d[22]),
    .c(al_a23f6f13),
    .o({al_52cd72b8,al_df3b43b5[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47384ade (
    .a(al_57dc9b0c[23]),
    .b(al_a5e9c08d[23]),
    .c(al_52cd72b8),
    .o({al_a35c5ad0,al_df3b43b5[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ffe133ad (
    .a(al_57dc9b0c[24]),
    .b(al_a5e9c08d[24]),
    .c(al_a35c5ad0),
    .o({al_bf78ad38,al_df3b43b5[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7fd6a45b (
    .a(al_57dc9b0c[25]),
    .b(al_a5e9c08d[25]),
    .c(al_bf78ad38),
    .o({al_f71c0797,al_df3b43b5[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3cb3fe3a (
    .a(al_57dc9b0c[26]),
    .b(al_a5e9c08d[26]),
    .c(al_f71c0797),
    .o({al_2d1a2942,al_df3b43b5[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_31e47287 (
    .a(al_57dc9b0c[0]),
    .b(al_a5e9c08d[0]),
    .c(al_bb31a1fd),
    .o({al_52f7b6db,al_df3b43b5[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a92c2cbc (
    .a(al_57dc9b0c[27]),
    .b(al_a5e9c08d[27]),
    .c(al_2d1a2942),
    .o({al_c045eda5,al_df3b43b5[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_43b69587 (
    .a(al_57dc9b0c[28]),
    .b(al_a5e9c08d[28]),
    .c(al_c045eda5),
    .o({al_892befbc,al_df3b43b5[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3dbc1cd (
    .a(al_57dc9b0c[29]),
    .b(al_a5e9c08d[29]),
    .c(al_892befbc),
    .o({al_19974a3,al_df3b43b5[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_da986575 (
    .a(al_57dc9b0c[30]),
    .b(al_a5e9c08d[30]),
    .c(al_19974a3),
    .o({al_634f8236,al_df3b43b5[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb5c7052 (
    .a(al_57dc9b0c[31]),
    .b(al_a5e9c08d[31]),
    .c(al_634f8236),
    .o({al_f607f1c2,al_df3b43b5[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d9f08d8 (
    .a(1'b0),
    .b(1'b1),
    .c(al_f607f1c2),
    .o({open_n129,al_42f85898}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff6125b (
    .a(al_57dc9b0c[1]),
    .b(al_a5e9c08d[1]),
    .c(al_52f7b6db),
    .o({al_a8fa8fea,al_df3b43b5[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_243d0ee5 (
    .a(al_57dc9b0c[2]),
    .b(al_a5e9c08d[2]),
    .c(al_a8fa8fea),
    .o({al_b2ffd084,al_df3b43b5[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a03b8532 (
    .a(al_57dc9b0c[3]),
    .b(al_a5e9c08d[3]),
    .c(al_b2ffd084),
    .o({al_b701d480,al_df3b43b5[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9cd7aa82 (
    .a(al_57dc9b0c[4]),
    .b(al_a5e9c08d[4]),
    .c(al_b701d480),
    .o({al_97262af6,al_df3b43b5[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a4b8a164 (
    .a(al_57dc9b0c[5]),
    .b(al_a5e9c08d[5]),
    .c(al_97262af6),
    .o({al_2a480b9e,al_df3b43b5[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9109a9ee (
    .a(al_57dc9b0c[6]),
    .b(al_a5e9c08d[6]),
    .c(al_2a480b9e),
    .o({al_d720b206,al_df3b43b5[6]}));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_57b13c7b (
    .a(al_dc0ce6da),
    .b(al_90a06cdf),
    .c(al_ecc3713),
    .d(al_4a1ebbca),
    .o(al_9535661e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_706d3730 (
    .a(al_b052c226[48]),
    .b(al_b052c226[49]),
    .c(al_b052c226[50]),
    .d(al_b052c226[51]),
    .e(al_b052c226[52]),
    .f(al_b052c226[53]),
    .o(al_3b37ef98));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_ea6046cb (
    .a(al_8691ef65),
    .b(al_b052c226[32]),
    .c(al_b052c226[33]),
    .d(al_b052c226[34]),
    .e(al_b052c226[35]),
    .o(al_ecc3713));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_cf2502f3 (
    .a(al_b052c226[44]),
    .b(al_b052c226[45]),
    .o(al_de5112e6));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_e64eb8e8 (
    .a(al_b052c226[46]),
    .b(al_b052c226[47]),
    .o(al_6c82a93e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_a2ff1fe9 (
    .a(al_de5112e6),
    .b(al_6c82a93e),
    .c(al_b052c226[40]),
    .d(al_b052c226[41]),
    .e(al_b052c226[42]),
    .f(al_b052c226[43]),
    .o(al_4a1ebbca));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_1fa7369f (
    .a(al_dc0ce6da),
    .b(al_90a06cdf),
    .c(al_ecc3713),
    .d(al_4a1ebbca),
    .e(al_b052c226[28]),
    .f(al_592f1b09[28]),
    .o(al_8c015879[28]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_86f0730c (
    .a(al_b052c226[56]),
    .b(al_b052c226[57]),
    .c(al_b052c226[58]),
    .d(al_b052c226[59]),
    .o(al_d63c55c7));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_102bacb1 (
    .a(al_3b37ef98),
    .b(al_d63c55c7),
    .c(al_b052c226[54]),
    .d(al_b052c226[55]),
    .o(al_dc0ce6da));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((~D*A))*~(E)*~(F)+~(B)*~(C)*~((~D*A))*E*~(F)+B*~(C)*~((~D*A))*E*~(F)+~(B)*~(C)*(~D*A)*E*~(F)+~(B)*~(C)*~((~D*A))*~(E)*F+B*~(C)*~((~D*A))*~(E)*F+~(B)*C*~((~D*A))*~(E)*F+~(B)*~(C)*(~D*A)*~(E)*F+B*~(C)*(~D*A)*~(E)*F+~(B)*~(C)*~((~D*A))*E*F+B*~(C)*~((~D*A))*E*F+~(B)*C*~((~D*A))*E*F+B*C*~((~D*A))*E*F+~(B)*~(C)*(~D*A)*E*F+B*~(C)*(~D*A)*E*F+~(B)*C*(~D*A)*E*F)"),
    .INIT(64'hff7f3f1f0f070301))
    al_c5c4bfa3 (
    .a(al_b052c226[28]),
    .b(al_b052c226[29]),
    .c(al_b052c226[30]),
    .d(al_592f1b09[28]),
    .e(al_592f1b09[29]),
    .f(al_592f1b09[30]),
    .o(al_7269924));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd4))
    al_fce89aa2 (
    .a(al_b052c226[31]),
    .b(al_592f1b09[31]),
    .c(al_7269924),
    .o(al_90a06cdf));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_231b6757 (
    .a(al_b052c226[36]),
    .b(al_b052c226[37]),
    .c(al_b052c226[38]),
    .d(al_b052c226[39]),
    .o(al_8691ef65));
  AL_MAP_LUT4 #(
    .EQN("~(D@B@(~C*A))"),
    .INIT(16'hc639))
    al_804bb09e (
    .a(al_b052c226[28]),
    .b(al_b052c226[29]),
    .c(al_592f1b09[28]),
    .d(al_592f1b09[29]),
    .o(al_54056c79));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E)*~((D*C*B*A))+~F*E*~((D*C*B*A))+~(~F)*E*(D*C*B*A)+~F*E*(D*C*B*A))"),
    .INIT(64'h7fffffff00008000))
    al_cc46c02a (
    .a(al_dc0ce6da),
    .b(al_90a06cdf),
    .c(al_ecc3713),
    .d(al_4a1ebbca),
    .e(al_54056c79),
    .f(al_592f1b09[29]),
    .o(al_8c015879[29]));
  AL_MAP_LUT6 #(
    .EQN("(F@C@(B*~((~D*A))*~(E)+~(B)*(~D*A)*~(E)+B*(~D*A)*~(E)+B*(~D*A)*E))"),
    .INIT(64'h0f87c3e1f0783c1e))
    al_1222e07c (
    .a(al_b052c226[28]),
    .b(al_b052c226[29]),
    .c(al_b052c226[30]),
    .d(al_592f1b09[28]),
    .e(al_592f1b09[29]),
    .f(al_592f1b09[30]),
    .o(al_828cf6c5[2]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E)*~((D*C*B*A))+F*E*~((D*C*B*A))+~(F)*E*(D*C*B*A)+F*E*(D*C*B*A))"),
    .INIT(64'hffff7fff80000000))
    al_f8267ca3 (
    .a(al_dc0ce6da),
    .b(al_90a06cdf),
    .c(al_ecc3713),
    .d(al_4a1ebbca),
    .e(al_828cf6c5[2]),
    .f(al_592f1b09[30]),
    .o(al_8c015879[30]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(C*B*A*~(E@D)))"),
    .INIT(64'h7fffff7f00000000))
    al_1a14712 (
    .a(al_dc0ce6da),
    .b(al_ecc3713),
    .c(al_4a1ebbca),
    .d(al_7269924),
    .e(al_b052c226[31]),
    .f(al_592f1b09[31]),
    .o(al_8c015879[31]));
  AL_DFF_X al_b824405e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44882eca[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f336c405[0]));
  AL_DFF_X al_629edd14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[27]));
  AL_DFF_X al_f4a37a2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[28]));
  AL_DFF_X al_8edfea8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[29]));
  AL_DFF_X al_78535658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[30]));
  AL_DFF_X al_206b9410 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[31]));
  AL_DFF_X al_cb054e86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[32]));
  AL_DFF_X al_ea1be463 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[33]));
  AL_DFF_X al_2829ee4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[34]));
  AL_DFF_X al_b2f1a406 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[35]));
  AL_DFF_X al_e90ca3b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[36]));
  AL_DFF_X al_ead04ad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[37]));
  AL_DFF_X al_e6d78dc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[38]));
  AL_DFF_X al_351c9015 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[39]));
  AL_DFF_X al_7597b4da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[40]));
  AL_DFF_X al_7affe042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[41]));
  AL_DFF_X al_1a2713ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[42]));
  AL_DFF_X al_c5e35689 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[43]));
  AL_DFF_X al_d986f01a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[44]));
  AL_DFF_X al_db244a97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[45]));
  AL_DFF_X al_86e0bf67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[46]));
  AL_DFF_X al_14043064 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[47]));
  AL_DFF_X al_4ac26836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[48]));
  AL_DFF_X al_94639f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[49]));
  AL_DFF_X al_d8b3455 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[50]));
  AL_DFF_X al_915db1b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[51]));
  AL_DFF_X al_664a0c46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[52]));
  AL_DFF_X al_54246cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[53]));
  AL_DFF_X al_1528e232 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[54]));
  AL_DFF_X al_26621aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[55]));
  AL_DFF_X al_4112dbd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[56]));
  AL_DFF_X al_f8aeace5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[57]));
  AL_DFF_X al_a739902b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[58]));
  AL_DFF_X al_7bca5b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[8]));
  AL_DFF_X al_95c635b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[9]));
  AL_DFF_X al_f828efc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[10]));
  AL_DFF_X al_91fdfa35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[11]));
  AL_DFF_X al_5a2b061 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[12]));
  AL_DFF_X al_a1e00e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[13]));
  AL_DFF_X al_5b84c1bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[14]));
  AL_DFF_X al_187c7814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[15]));
  AL_DFF_X al_1871d527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[16]));
  AL_DFF_X al_42ca7269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[17]));
  AL_DFF_X al_24e134af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[0]));
  AL_DFF_X al_29a5ac71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[18]));
  AL_DFF_X al_d5f7e29e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[19]));
  AL_DFF_X al_8a96d3e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[20]));
  AL_DFF_X al_240ad317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[21]));
  AL_DFF_X al_abd74ff6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[22]));
  AL_DFF_X al_55a527d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[23]));
  AL_DFF_X al_f479891a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[24]));
  AL_DFF_X al_afedc3fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[25]));
  AL_DFF_X al_53b5c590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[26]));
  AL_DFF_X al_c053b796 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[27]));
  AL_DFF_X al_141a1472 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[1]));
  AL_DFF_X al_e26e15e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[28]));
  AL_DFF_X al_dfa0cc31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[29]));
  AL_DFF_X al_8a901de9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[30]));
  AL_DFF_X al_7597602c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[31]));
  AL_DFF_X al_2aaa9264 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[2]));
  AL_DFF_X al_855d6b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[3]));
  AL_DFF_X al_1759d677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[4]));
  AL_DFF_X al_e3ab410d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[5]));
  AL_DFF_X al_1f370737 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[6]));
  AL_DFF_X al_90e5a34b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[7]));
  AL_DFF_X al_6004626e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9535661e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[0]));
  AL_DFF_X al_e60ff7a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[1]));
  AL_DFF_X al_a1b664a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[2]));
  AL_DFF_X al_7c1acbb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ffc2fb62 (
    .a(al_57ac52e7),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .o(al_2be1d9b7));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((~D*A))*~(E)*~(F)+~(B)*~(C)*~((~D*A))*E*~(F)+B*~(C)*~((~D*A))*E*~(F)+~(B)*~(C)*(~D*A)*E*~(F)+~(B)*~(C)*~((~D*A))*~(E)*F+B*~(C)*~((~D*A))*~(E)*F+~(B)*C*~((~D*A))*~(E)*F+~(B)*~(C)*(~D*A)*~(E)*F+B*~(C)*(~D*A)*~(E)*F+~(B)*~(C)*~((~D*A))*E*F+B*~(C)*~((~D*A))*E*F+~(B)*C*~((~D*A))*E*F+B*C*~((~D*A))*E*F+~(B)*~(C)*(~D*A)*E*F+B*~(C)*(~D*A)*E*F+~(B)*C*(~D*A)*E*F)"),
    .INIT(64'hff7f3f1f0f070301))
    al_b5111bba (
    .a(al_28202fa7[27]),
    .b(al_28202fa7[28]),
    .c(al_28202fa7[29]),
    .d(al_1d4399b1[27]),
    .e(al_1d4399b1[28]),
    .f(al_1d4399b1[29]),
    .o(al_4f7fb1ad));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_b4a36fc3 (
    .a(al_cadea4c8),
    .b(al_28202fa7[32]),
    .c(al_28202fa7[35]),
    .d(al_28202fa7[37]),
    .e(al_28202fa7[38]),
    .o(al_203d257f));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_31e32617 (
    .a(al_28202fa7[56]),
    .b(al_28202fa7[57]),
    .o(al_ca8f2e4c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_fb49539c (
    .a(al_ca8f2e4c),
    .b(al_28202fa7[48]),
    .c(al_28202fa7[51]),
    .d(al_28202fa7[53]),
    .e(al_28202fa7[54]),
    .f(al_28202fa7[58]),
    .o(al_ed33bb97));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_1ad31b56 (
    .a(al_57ac52e7),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .e(al_28202fa7[27]),
    .f(al_1d4399b1[27]),
    .o(al_7a8c14f1[27]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbf2f0b02))
    al_4b55cad3 (
    .a(al_4f7fb1ad),
    .b(al_28202fa7[30]),
    .c(al_28202fa7[31]),
    .d(al_1d4399b1[30]),
    .e(al_1d4399b1[31]),
    .o(al_57ac52e7));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_fc152134 (
    .a(al_28202fa7[49]),
    .b(al_28202fa7[50]),
    .c(al_28202fa7[52]),
    .d(al_28202fa7[55]),
    .o(al_1e591849));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_fcfa038 (
    .a(al_28202fa7[36]),
    .b(al_28202fa7[39]),
    .c(al_28202fa7[40]),
    .d(al_28202fa7[43]),
    .o(al_e40698dd));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_da80ede8 (
    .a(al_1e591849),
    .b(al_e40698dd),
    .c(al_28202fa7[33]),
    .d(al_28202fa7[34]),
    .e(al_28202fa7[45]),
    .f(al_28202fa7[46]),
    .o(al_552d5319));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_412eaacf (
    .a(al_28202fa7[41]),
    .b(al_28202fa7[42]),
    .c(al_28202fa7[44]),
    .d(al_28202fa7[47]),
    .o(al_cadea4c8));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b9028d97 (
    .a(al_28202fa7[27]),
    .b(al_1d4399b1[27]),
    .o(al_82784f18));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e7e1a754 (
    .a(al_82784f18),
    .b(al_28202fa7[28]),
    .o(al_2281381d));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_2a00686 (
    .a(al_57ac52e7),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .e(al_2281381d),
    .f(al_1d4399b1[28]),
    .o(al_7a8c14f1[28]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    .INIT(16'h781e))
    al_2e5ee078 (
    .a(al_82784f18),
    .b(al_28202fa7[28]),
    .c(al_28202fa7[29]),
    .d(al_1d4399b1[28]),
    .o(al_2f03a26));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_5c102dbd (
    .a(al_57ac52e7),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .e(al_2f03a26),
    .f(al_1d4399b1[29]),
    .o(al_7a8c14f1[29]));
  AL_MAP_LUT6 #(
    .EQN("(D@(~(A)*~(B)*~(C)*~(E)*~(F)+~(A)*~(B)*~(C)*E*~(F)+A*~(B)*~(C)*E*~(F)+~(A)*B*~(C)*E*~(F)+~(A)*~(B)*~(C)*~(E)*F+A*~(B)*~(C)*~(E)*F+~(A)*B*~(C)*~(E)*F+A*B*~(C)*~(E)*F+~(A)*~(B)*C*~(E)*F+~(A)*~(B)*~(C)*E*F+A*~(B)*~(C)*E*F+~(A)*B*~(C)*E*F+A*B*~(C)*E*F+~(A)*~(B)*C*E*F+A*~(B)*C*E*F+~(A)*B*C*E*F))"),
    .INIT(64'h807fe01ff807fe01))
    al_b1151c99 (
    .a(al_82784f18),
    .b(al_28202fa7[28]),
    .c(al_28202fa7[29]),
    .d(al_28202fa7[30]),
    .e(al_1d4399b1[28]),
    .f(al_1d4399b1[29]),
    .o(al_6f00a1da));
  AL_MAP_LUT6 #(
    .EQN("(F@(~E*D*C*B*A))"),
    .INIT(64'hffff7fff00008000))
    al_af9fc655 (
    .a(al_57ac52e7),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .e(al_6f00a1da),
    .f(al_1d4399b1[30]),
    .o(al_7a8c14f1[30]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*B*C)"),
    .INIT(8'h4d))
    al_d3f46475 (
    .a(al_4f7fb1ad),
    .b(al_28202fa7[30]),
    .c(al_1d4399b1[30]),
    .o(al_f96974bd));
  AL_MAP_LUT6 #(
    .EQN("(F*~(D*C*B*(E@A)))"),
    .INIT(64'hbfff7fff00000000))
    al_7d8fa9e8 (
    .a(al_f96974bd),
    .b(al_552d5319),
    .c(al_203d257f),
    .d(al_ed33bb97),
    .e(al_28202fa7[31]),
    .f(al_1d4399b1[31]),
    .o(al_7a8c14f1[31]));
  AL_DFF_X al_c1b05d22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f336c405[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f23786d8[0]));
  AL_DFF_X al_16c9a7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[26]));
  AL_DFF_X al_74f6e083 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[27]));
  AL_DFF_X al_4e512437 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[28]));
  AL_DFF_X al_db10517f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[29]));
  AL_DFF_X al_c6183e37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[30]));
  AL_DFF_X al_4f2a5e19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[31]));
  AL_DFF_X al_2d3ce6cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[32]));
  AL_DFF_X al_88919bdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[33]));
  AL_DFF_X al_90109587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[34]));
  AL_DFF_X al_74d431c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[35]));
  AL_DFF_X al_2d99e7e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[36]));
  AL_DFF_X al_9b5e8323 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[37]));
  AL_DFF_X al_edfc91bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[38]));
  AL_DFF_X al_4ec3bd0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[39]));
  AL_DFF_X al_bea2a272 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[40]));
  AL_DFF_X al_4411ed5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[41]));
  AL_DFF_X al_85376b89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[42]));
  AL_DFF_X al_e6428e2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[43]));
  AL_DFF_X al_6e673a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[44]));
  AL_DFF_X al_b321bddc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[45]));
  AL_DFF_X al_a33a4af3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[46]));
  AL_DFF_X al_23d2a568 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[47]));
  AL_DFF_X al_1515111b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[48]));
  AL_DFF_X al_a8fbb28c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[49]));
  AL_DFF_X al_80c553a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[50]));
  AL_DFF_X al_1d749880 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[51]));
  AL_DFF_X al_607edc2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[52]));
  AL_DFF_X al_4cd3ae3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[53]));
  AL_DFF_X al_714444c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[54]));
  AL_DFF_X al_34814d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[55]));
  AL_DFF_X al_df74699a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[56]));
  AL_DFF_X al_a8fd7641 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[57]));
  AL_DFF_X al_30045b86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[8]));
  AL_DFF_X al_30c4a0cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[9]));
  AL_DFF_X al_ccd54ad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[10]));
  AL_DFF_X al_a346acb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[11]));
  AL_DFF_X al_52728c4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[12]));
  AL_DFF_X al_defcd91c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[13]));
  AL_DFF_X al_f58d7987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[14]));
  AL_DFF_X al_d26f4b8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[15]));
  AL_DFF_X al_11702fae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[16]));
  AL_DFF_X al_bd8c811d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[17]));
  AL_DFF_X al_29600c3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[0]));
  AL_DFF_X al_50b9e82e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[18]));
  AL_DFF_X al_44a652d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[19]));
  AL_DFF_X al_e1cfc4d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[20]));
  AL_DFF_X al_eb87b308 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[21]));
  AL_DFF_X al_35bd6a86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[22]));
  AL_DFF_X al_d6a4c3fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[23]));
  AL_DFF_X al_fc6f72b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[24]));
  AL_DFF_X al_a2cd993d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[25]));
  AL_DFF_X al_7c4cbd84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[26]));
  AL_DFF_X al_8ed23af2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[27]));
  AL_DFF_X al_8b3164c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[1]));
  AL_DFF_X al_fe47a994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[28]));
  AL_DFF_X al_71230d17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[29]));
  AL_DFF_X al_3bc55982 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[30]));
  AL_DFF_X al_9836f82f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[31]));
  AL_DFF_X al_9a3602d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[2]));
  AL_DFF_X al_e50f91fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[3]));
  AL_DFF_X al_f4e16c6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[4]));
  AL_DFF_X al_e188fed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[5]));
  AL_DFF_X al_1c2aa46a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[6]));
  AL_DFF_X al_dd3656c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[7]));
  AL_DFF_X al_dc4ef4ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2be1d9b7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[0]));
  AL_DFF_X al_8d8268f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[1]));
  AL_DFF_X al_14b0d265 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[2]));
  AL_DFF_X al_46ba5fed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[3]));
  AL_DFF_X al_aef1e997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8605901e (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .o(al_f3cdefe2));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_fa102b68 (
    .a(1'b0),
    .o({al_5f980ce9,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec0ccb55 (
    .a(al_1b3e91c5[26]),
    .b(al_68bb3ebd[26]),
    .c(al_5f980ce9),
    .o({al_a2de35e1,al_d01f30c3[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b5f4de94 (
    .a(al_1b3e91c5[27]),
    .b(al_68bb3ebd[27]),
    .c(al_a2de35e1),
    .o({al_4ba9ed11,al_d01f30c3[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c4391072 (
    .a(al_1b3e91c5[28]),
    .b(al_68bb3ebd[28]),
    .c(al_4ba9ed11),
    .o({al_cacb9d80,al_d01f30c3[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a0d30c4 (
    .a(al_1b3e91c5[29]),
    .b(al_68bb3ebd[29]),
    .c(al_cacb9d80),
    .o({al_1bad0a7d,al_d01f30c3[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8f3c8801 (
    .a(al_1b3e91c5[30]),
    .b(al_68bb3ebd[30]),
    .c(al_1bad0a7d),
    .o({al_58234d6b,al_d01f30c3[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a1bbffc8 (
    .a(al_1b3e91c5[31]),
    .b(al_68bb3ebd[31]),
    .c(al_58234d6b),
    .o({al_c5f2b310,al_d01f30c3[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1d7430b (
    .c(al_c5f2b310),
    .o({open_n135,al_d01f30c3[6]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_40358306 (
    .a(al_68bb3ebd[46]),
    .b(al_68bb3ebd[47]),
    .c(al_68bb3ebd[48]),
    .d(al_68bb3ebd[49]),
    .e(al_68bb3ebd[50]),
    .f(al_68bb3ebd[51]),
    .o(al_477c87));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_312525b2 (
    .a(al_68bb3ebd[36]),
    .b(al_68bb3ebd[37]),
    .c(al_68bb3ebd[38]),
    .d(al_68bb3ebd[39]),
    .o(al_b8df04a0));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_629f3954 (
    .a(al_cb5c1242),
    .b(al_b8df04a0),
    .c(al_68bb3ebd[34]),
    .d(al_68bb3ebd[35]),
    .e(al_68bb3ebd[40]),
    .f(al_68bb3ebd[41]),
    .o(al_93714d98));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_d37cedfd (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[26]),
    .d(al_d01f30c3[0]),
    .o(al_7d7cdb8e[26]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_5c8b85ce (
    .a(al_68bb3ebd[54]),
    .b(al_68bb3ebd[55]),
    .c(al_68bb3ebd[56]),
    .d(al_68bb3ebd[57]),
    .o(al_b103a97e));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_e82a0a45 (
    .a(al_68bb3ebd[32]),
    .b(al_68bb3ebd[33]),
    .c(al_d01f30c3[6]),
    .o(al_d405f4db));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_9a754097 (
    .a(al_477c87),
    .b(al_b103a97e),
    .c(al_d405f4db),
    .d(al_68bb3ebd[52]),
    .e(al_68bb3ebd[53]),
    .o(al_59bc69f9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_c630ac94 (
    .a(al_68bb3ebd[42]),
    .b(al_68bb3ebd[43]),
    .c(al_68bb3ebd[44]),
    .d(al_68bb3ebd[45]),
    .o(al_cb5c1242));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_7147c201 (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[27]),
    .d(al_d01f30c3[1]),
    .o(al_7d7cdb8e[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_188ceff (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[28]),
    .d(al_d01f30c3[2]),
    .o(al_7d7cdb8e[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_4e202a7a (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[29]),
    .d(al_d01f30c3[3]),
    .o(al_7d7cdb8e[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_32724b32 (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[30]),
    .d(al_d01f30c3[4]),
    .o(al_7d7cdb8e[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_78d63c10 (
    .a(al_59bc69f9),
    .b(al_93714d98),
    .c(al_1b3e91c5[31]),
    .d(al_d01f30c3[5]),
    .o(al_7d7cdb8e[31]));
  AL_DFF_X al_4e46745 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f23786d8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6e4d5f5f[0]));
  AL_DFF_X al_2c1c2b5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[25]));
  AL_DFF_X al_4801a8af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[26]));
  AL_DFF_X al_d0e21fb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[27]));
  AL_DFF_X al_d9db21a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[28]));
  AL_DFF_X al_ef12853f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[29]));
  AL_DFF_X al_bd29404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[30]));
  AL_DFF_X al_4d4abdfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[31]));
  AL_DFF_X al_fc1d6c08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[32]));
  AL_DFF_X al_ec0464b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[33]));
  AL_DFF_X al_a8789532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[34]));
  AL_DFF_X al_9c63114d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[35]));
  AL_DFF_X al_b9bf9d2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[36]));
  AL_DFF_X al_28a3e61e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[37]));
  AL_DFF_X al_ba3c61a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[38]));
  AL_DFF_X al_bceccfbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[39]));
  AL_DFF_X al_17c2ceeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[40]));
  AL_DFF_X al_d7332f93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[41]));
  AL_DFF_X al_dcf8608d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[42]));
  AL_DFF_X al_f574ae6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[43]));
  AL_DFF_X al_e90f82f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[44]));
  AL_DFF_X al_7fd1efb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[45]));
  AL_DFF_X al_faff71e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[46]));
  AL_DFF_X al_fcc61d29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[47]));
  AL_DFF_X al_d46b7da7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[48]));
  AL_DFF_X al_ee2311bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[49]));
  AL_DFF_X al_3b6761cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[50]));
  AL_DFF_X al_c6092adb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[51]));
  AL_DFF_X al_6b43d194 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[52]));
  AL_DFF_X al_ea5f28a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[53]));
  AL_DFF_X al_12538005 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[54]));
  AL_DFF_X al_1fae0736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[55]));
  AL_DFF_X al_451ffb8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[56]));
  AL_DFF_X al_d1ea0b4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[8]));
  AL_DFF_X al_6566d01e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[9]));
  AL_DFF_X al_9cc2148c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[10]));
  AL_DFF_X al_1adf66fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[11]));
  AL_DFF_X al_d6ee48a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[12]));
  AL_DFF_X al_d65ad79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[13]));
  AL_DFF_X al_c8b5ec82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[14]));
  AL_DFF_X al_119001 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[15]));
  AL_DFF_X al_635da4e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[16]));
  AL_DFF_X al_b3bd2fea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[17]));
  AL_DFF_X al_b8837cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[0]));
  AL_DFF_X al_1f79729a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[18]));
  AL_DFF_X al_87ed3178 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[19]));
  AL_DFF_X al_20c2fb5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[20]));
  AL_DFF_X al_b6e21ad6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[21]));
  AL_DFF_X al_d8bd7831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[22]));
  AL_DFF_X al_4d4ec29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[23]));
  AL_DFF_X al_eb3b77cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[24]));
  AL_DFF_X al_b366953f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[25]));
  AL_DFF_X al_a335f641 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[26]));
  AL_DFF_X al_88b23d06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[27]));
  AL_DFF_X al_2205221c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[1]));
  AL_DFF_X al_63814eb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[28]));
  AL_DFF_X al_e5676122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[29]));
  AL_DFF_X al_c231fa47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[30]));
  AL_DFF_X al_173f8e20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[31]));
  AL_DFF_X al_f82771e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[2]));
  AL_DFF_X al_49d9b260 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[3]));
  AL_DFF_X al_1f30d5c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[4]));
  AL_DFF_X al_a9722f97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[5]));
  AL_DFF_X al_4a6c2985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[6]));
  AL_DFF_X al_f7736fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[7]));
  AL_DFF_X al_ca9d3a14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3cdefe2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[0]));
  AL_DFF_X al_5cec555d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[1]));
  AL_DFF_X al_f35bc942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[2]));
  AL_DFF_X al_af6b3c25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[3]));
  AL_DFF_X al_2e20cd82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[4]));
  AL_DFF_X al_b7748714 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fd4ffc73 (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .o(al_4de4f552));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ed11b73e (
    .a(1'b0),
    .o({al_25f6edd0,open_n138}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68fbbe18 (
    .a(al_15503509[25]),
    .b(al_f2a9de02[25]),
    .c(al_25f6edd0),
    .o({al_4b9b0b4,al_f3dd9213[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40bfb914 (
    .a(al_15503509[26]),
    .b(al_f2a9de02[26]),
    .c(al_4b9b0b4),
    .o({al_4ecce1a8,al_f3dd9213[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_15108eaf (
    .a(al_15503509[27]),
    .b(al_f2a9de02[27]),
    .c(al_4ecce1a8),
    .o({al_a74a382d,al_f3dd9213[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2316cbde (
    .a(al_15503509[28]),
    .b(al_f2a9de02[28]),
    .c(al_a74a382d),
    .o({al_fa0c3c8b,al_f3dd9213[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_750b81ba (
    .a(al_15503509[29]),
    .b(al_f2a9de02[29]),
    .c(al_fa0c3c8b),
    .o({al_67ed9c11,al_f3dd9213[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27b5d17c (
    .a(al_15503509[30]),
    .b(al_f2a9de02[30]),
    .c(al_67ed9c11),
    .o({al_f563230a,al_f3dd9213[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9de1adb (
    .a(al_15503509[31]),
    .b(al_f2a9de02[31]),
    .c(al_f563230a),
    .o({al_c539d3e8,al_f3dd9213[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ecff783b (
    .c(al_c539d3e8),
    .o({open_n141,al_f3dd9213[7]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_8fc9c265 (
    .a(al_f2a9de02[34]),
    .b(al_f2a9de02[35]),
    .c(al_f2a9de02[36]),
    .d(al_f2a9de02[37]),
    .e(al_f2a9de02[38]),
    .f(al_f2a9de02[39]),
    .o(al_79960e7c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_ffd23aee (
    .a(al_631391e1),
    .b(al_126d5412),
    .c(al_f2a9de02[46]),
    .d(al_f2a9de02[47]),
    .e(al_f2a9de02[52]),
    .f(al_f2a9de02[53]),
    .o(al_7c9dcdbf));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_a7660868 (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[25]),
    .d(al_f3dd9213[0]),
    .o(al_78306f09[25]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_ef108187 (
    .a(al_f2a9de02[42]),
    .b(al_f2a9de02[43]),
    .c(al_f2a9de02[44]),
    .d(al_f2a9de02[45]),
    .o(al_a9fdceb9));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_3458a018 (
    .a(al_79960e7c),
    .b(al_a9fdceb9),
    .c(al_f2a9de02[32]),
    .d(al_f2a9de02[33]),
    .e(al_f2a9de02[40]),
    .f(al_f2a9de02[41]),
    .o(al_c9a744c1));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6dc5abdc (
    .a(al_f2a9de02[54]),
    .b(al_f2a9de02[55]),
    .c(al_f2a9de02[56]),
    .d(al_f3dd9213[7]),
    .o(al_631391e1));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_901e07bd (
    .a(al_f2a9de02[48]),
    .b(al_f2a9de02[49]),
    .c(al_f2a9de02[50]),
    .d(al_f2a9de02[51]),
    .o(al_126d5412));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ee0ec1c (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[26]),
    .d(al_f3dd9213[1]),
    .o(al_78306f09[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_ee73087c (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[27]),
    .d(al_f3dd9213[2]),
    .o(al_78306f09[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_42a9db3d (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[28]),
    .d(al_f3dd9213[3]),
    .o(al_78306f09[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_a11411b (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[29]),
    .d(al_f3dd9213[4]),
    .o(al_78306f09[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_cee49f18 (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[30]),
    .d(al_f3dd9213[5]),
    .o(al_78306f09[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9aa0eda8 (
    .a(al_c9a744c1),
    .b(al_7c9dcdbf),
    .c(al_15503509[31]),
    .d(al_f3dd9213[6]),
    .o(al_78306f09[31]));
  AL_DFF_X al_54bb73dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6e4d5f5f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d255f877[0]));
  AL_DFF_X al_cf7645d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[24]));
  AL_DFF_X al_3fefb87b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[25]));
  AL_DFF_X al_1a9ac779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[26]));
  AL_DFF_X al_36aa0f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[27]));
  AL_DFF_X al_925290f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[28]));
  AL_DFF_X al_b9345772 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[29]));
  AL_DFF_X al_f7413fa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[30]));
  AL_DFF_X al_545fe956 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[31]));
  AL_DFF_X al_c4167b1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[32]));
  AL_DFF_X al_4963703f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[33]));
  AL_DFF_X al_2eaa9255 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[34]));
  AL_DFF_X al_5cd3f66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[35]));
  AL_DFF_X al_2770fff1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[36]));
  AL_DFF_X al_2fb88ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[37]));
  AL_DFF_X al_33188a38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[38]));
  AL_DFF_X al_518187d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[39]));
  AL_DFF_X al_5086df15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[40]));
  AL_DFF_X al_8f4fd57c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[41]));
  AL_DFF_X al_f17c1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[42]));
  AL_DFF_X al_788e73ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[43]));
  AL_DFF_X al_fac2367e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[44]));
  AL_DFF_X al_5525468a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[45]));
  AL_DFF_X al_205e1075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[46]));
  AL_DFF_X al_f657423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[47]));
  AL_DFF_X al_d1be2a7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[48]));
  AL_DFF_X al_40063a27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[49]));
  AL_DFF_X al_6928b682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[50]));
  AL_DFF_X al_1751be99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[51]));
  AL_DFF_X al_f1fd591b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[52]));
  AL_DFF_X al_ad7b5bfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[53]));
  AL_DFF_X al_b4fa4244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[54]));
  AL_DFF_X al_be11be3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[55]));
  AL_DFF_X al_1afa1258 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[8]));
  AL_DFF_X al_71a16da7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[9]));
  AL_DFF_X al_7d507b3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[10]));
  AL_DFF_X al_59921bf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[11]));
  AL_DFF_X al_661a65b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[12]));
  AL_DFF_X al_280330c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[13]));
  AL_DFF_X al_ba352714 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[14]));
  AL_DFF_X al_5c43f732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[15]));
  AL_DFF_X al_a35b6858 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[16]));
  AL_DFF_X al_cbf371c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[17]));
  AL_DFF_X al_77c3e7d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[0]));
  AL_DFF_X al_fa109aec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[18]));
  AL_DFF_X al_eca2af20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[19]));
  AL_DFF_X al_392585f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[20]));
  AL_DFF_X al_3ca470de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[21]));
  AL_DFF_X al_a219939f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[22]));
  AL_DFF_X al_a8ef659a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[23]));
  AL_DFF_X al_df040b95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[24]));
  AL_DFF_X al_643f4509 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[25]));
  AL_DFF_X al_7f4c7397 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[26]));
  AL_DFF_X al_d3b08ec4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[27]));
  AL_DFF_X al_fb19511f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[1]));
  AL_DFF_X al_da75108b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[28]));
  AL_DFF_X al_afc07418 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[29]));
  AL_DFF_X al_dbb3cd36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[30]));
  AL_DFF_X al_afbfc9f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[31]));
  AL_DFF_X al_f84305c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[2]));
  AL_DFF_X al_c5253883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[3]));
  AL_DFF_X al_3061a46b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[4]));
  AL_DFF_X al_a219d325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[5]));
  AL_DFF_X al_a66cb14f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[6]));
  AL_DFF_X al_826b2a64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[7]));
  AL_DFF_X al_31602fe8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4de4f552),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[0]));
  AL_DFF_X al_e39fd14b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[1]));
  AL_DFF_X al_bfef8c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[2]));
  AL_DFF_X al_c6ca6313 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[3]));
  AL_DFF_X al_c521ec6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[4]));
  AL_DFF_X al_aaaf72da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[5]));
  AL_DFF_X al_525dc2be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7175fe4a (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .o(al_1fc14639));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_51515bf (
    .a(1'b0),
    .o({al_753472e,open_n144}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f461f14 (
    .a(al_59bef53b[24]),
    .b(al_5206392b[24]),
    .c(al_753472e),
    .o({al_15e33bf2,al_727f921[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52bf100a (
    .a(al_59bef53b[25]),
    .b(al_5206392b[25]),
    .c(al_15e33bf2),
    .o({al_64c930a8,al_727f921[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6af7a3fe (
    .a(al_59bef53b[26]),
    .b(al_5206392b[26]),
    .c(al_64c930a8),
    .o({al_6ff407e,al_727f921[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_500a11b2 (
    .a(al_59bef53b[27]),
    .b(al_5206392b[27]),
    .c(al_6ff407e),
    .o({al_ff0e3144,al_727f921[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14355756 (
    .a(al_59bef53b[28]),
    .b(al_5206392b[28]),
    .c(al_ff0e3144),
    .o({al_f8599920,al_727f921[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_81bb53eb (
    .a(al_59bef53b[29]),
    .b(al_5206392b[29]),
    .c(al_f8599920),
    .o({al_b9af15ec,al_727f921[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c05631a2 (
    .a(al_59bef53b[30]),
    .b(al_5206392b[30]),
    .c(al_b9af15ec),
    .o({al_47c20a17,al_727f921[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9f255840 (
    .a(al_59bef53b[31]),
    .b(al_5206392b[31]),
    .c(al_47c20a17),
    .o({al_f5506553,al_727f921[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b39fd4e (
    .c(al_f5506553),
    .o({open_n147,al_727f921[8]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_dac50b62 (
    .a(al_5206392b[44]),
    .b(al_5206392b[45]),
    .c(al_5206392b[46]),
    .d(al_5206392b[47]),
    .e(al_5206392b[48]),
    .f(al_5206392b[49]),
    .o(al_a989c55e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_fb8ecff (
    .a(al_682ed5c4),
    .b(al_75a022),
    .c(al_5206392b[32]),
    .d(al_5206392b[33]),
    .e(al_5206392b[38]),
    .f(al_5206392b[39]),
    .o(al_81b3dbd9));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_60299857 (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[24]),
    .d(al_727f921[0]),
    .o(al_601b9c02[24]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_66c518e5 (
    .a(al_5206392b[52]),
    .b(al_5206392b[53]),
    .c(al_5206392b[54]),
    .d(al_5206392b[55]),
    .o(al_6dfedbe6));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_bd78d9af (
    .a(al_a989c55e),
    .b(al_6dfedbe6),
    .c(al_5206392b[50]),
    .d(al_5206392b[51]),
    .e(al_727f921[8]),
    .o(al_cce5b1fa));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_196a3474 (
    .a(al_5206392b[40]),
    .b(al_5206392b[41]),
    .c(al_5206392b[42]),
    .d(al_5206392b[43]),
    .o(al_682ed5c4));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6ab26684 (
    .a(al_5206392b[34]),
    .b(al_5206392b[35]),
    .c(al_5206392b[36]),
    .d(al_5206392b[37]),
    .o(al_75a022));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_f1ad9c4d (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[25]),
    .d(al_727f921[1]),
    .o(al_601b9c02[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_8522c1ef (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[26]),
    .d(al_727f921[2]),
    .o(al_601b9c02[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_c204cd0b (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[27]),
    .d(al_727f921[3]),
    .o(al_601b9c02[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_8565d196 (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[28]),
    .d(al_727f921[4]),
    .o(al_601b9c02[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_81935c6c (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[29]),
    .d(al_727f921[5]),
    .o(al_601b9c02[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_3d9f7478 (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[30]),
    .d(al_727f921[6]),
    .o(al_601b9c02[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_1f6007b8 (
    .a(al_cce5b1fa),
    .b(al_81b3dbd9),
    .c(al_59bef53b[31]),
    .d(al_727f921[7]),
    .o(al_601b9c02[31]));
  AL_DFF_X al_50e2d110 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d255f877[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30922aac[0]));
  AL_DFF_X al_31b6bc1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[23]));
  AL_DFF_X al_ed18db8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[24]));
  AL_DFF_X al_8a55ce2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[25]));
  AL_DFF_X al_61eaab3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[26]));
  AL_DFF_X al_29dc2cee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[27]));
  AL_DFF_X al_4ddc6ff4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[28]));
  AL_DFF_X al_10abbbc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[29]));
  AL_DFF_X al_9ae5bc94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[30]));
  AL_DFF_X al_8638d5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[31]));
  AL_DFF_X al_1154c404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[32]));
  AL_DFF_X al_f175541c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[33]));
  AL_DFF_X al_ec4f05a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[34]));
  AL_DFF_X al_ba6450cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[35]));
  AL_DFF_X al_2fa9f35e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[36]));
  AL_DFF_X al_3c9f056b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[37]));
  AL_DFF_X al_7b24af23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[38]));
  AL_DFF_X al_32bd1ac9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[39]));
  AL_DFF_X al_63d46252 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[40]));
  AL_DFF_X al_2434deaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[41]));
  AL_DFF_X al_28bbd23c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[42]));
  AL_DFF_X al_59d21a36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[43]));
  AL_DFF_X al_73de7de6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[44]));
  AL_DFF_X al_8def737f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[45]));
  AL_DFF_X al_5b0c2532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[46]));
  AL_DFF_X al_b8f8c880 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[47]));
  AL_DFF_X al_68223dba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[48]));
  AL_DFF_X al_624dac5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[49]));
  AL_DFF_X al_6b64e9c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[50]));
  AL_DFF_X al_8646f558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[51]));
  AL_DFF_X al_f539862f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[52]));
  AL_DFF_X al_951f469b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[53]));
  AL_DFF_X al_9031070f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[54]));
  AL_DFF_X al_dad62689 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[8]));
  AL_DFF_X al_4310eebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[9]));
  AL_DFF_X al_f566a5f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[10]));
  AL_DFF_X al_cbd3310b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[11]));
  AL_DFF_X al_5c978668 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[12]));
  AL_DFF_X al_b985e5b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[13]));
  AL_DFF_X al_1afa10a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[14]));
  AL_DFF_X al_fd28eb9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[15]));
  AL_DFF_X al_dbd7a2ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[16]));
  AL_DFF_X al_dc972ff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[17]));
  AL_DFF_X al_bbfb8607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[0]));
  AL_DFF_X al_340c32b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[18]));
  AL_DFF_X al_8e8fc704 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[19]));
  AL_DFF_X al_84ecb6aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[20]));
  AL_DFF_X al_6d41d36b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[21]));
  AL_DFF_X al_9792b3e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[22]));
  AL_DFF_X al_dfa0f87b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[23]));
  AL_DFF_X al_19ddb72a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[24]));
  AL_DFF_X al_625a9cbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[25]));
  AL_DFF_X al_f99ef2df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[26]));
  AL_DFF_X al_285865e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[27]));
  AL_DFF_X al_fe94433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[1]));
  AL_DFF_X al_cdef0355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[28]));
  AL_DFF_X al_506385c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[29]));
  AL_DFF_X al_e2766b77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[30]));
  AL_DFF_X al_de10ad32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[31]));
  AL_DFF_X al_90d2e951 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[2]));
  AL_DFF_X al_7986e6a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[3]));
  AL_DFF_X al_2f49a850 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[4]));
  AL_DFF_X al_1aa8b256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[5]));
  AL_DFF_X al_7582bb2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[6]));
  AL_DFF_X al_fbe03a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[7]));
  AL_DFF_X al_640a9d37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1fc14639),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[0]));
  AL_DFF_X al_6dfb03fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[1]));
  AL_DFF_X al_af6b473c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[2]));
  AL_DFF_X al_b7fee3ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[3]));
  AL_DFF_X al_a36ede7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[4]));
  AL_DFF_X al_26c44c89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[5]));
  AL_DFF_X al_6035cc5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[6]));
  AL_DFF_X al_69c1108d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_9f3aec89 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .o(al_d150e9d));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ed682aab (
    .a(1'b0),
    .o({al_d1df1e3c,open_n150}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9cb4768 (
    .a(al_f7a9a92b[23]),
    .b(al_d6cb04b6[23]),
    .c(al_d1df1e3c),
    .o({al_c46bddb5,al_96e7074d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_20eb07d7 (
    .a(al_f7a9a92b[24]),
    .b(al_d6cb04b6[24]),
    .c(al_c46bddb5),
    .o({al_24bfc94c,al_96e7074d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92c2cc99 (
    .a(al_f7a9a92b[25]),
    .b(al_d6cb04b6[25]),
    .c(al_24bfc94c),
    .o({al_92dd4899,al_96e7074d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a2cf30a9 (
    .a(al_f7a9a92b[26]),
    .b(al_d6cb04b6[26]),
    .c(al_92dd4899),
    .o({al_79a8092a,al_96e7074d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7572e88 (
    .a(al_f7a9a92b[27]),
    .b(al_d6cb04b6[27]),
    .c(al_79a8092a),
    .o({al_7e098907,al_96e7074d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a1084916 (
    .a(al_f7a9a92b[28]),
    .b(al_d6cb04b6[28]),
    .c(al_7e098907),
    .o({al_ad4f86b8,al_96e7074d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa6bd7bd (
    .a(al_f7a9a92b[29]),
    .b(al_d6cb04b6[29]),
    .c(al_ad4f86b8),
    .o({al_a5ca0ead,al_96e7074d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59e1a944 (
    .a(al_f7a9a92b[30]),
    .b(al_d6cb04b6[30]),
    .c(al_a5ca0ead),
    .o({al_ef88efba,al_96e7074d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f55eba23 (
    .a(al_f7a9a92b[31]),
    .b(al_d6cb04b6[31]),
    .c(al_ef88efba),
    .o({al_15966972,al_96e7074d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd4f3433 (
    .c(al_15966972),
    .o({open_n153,al_96e7074d[9]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b62ccded (
    .a(al_d6cb04b6[32]),
    .b(al_d6cb04b6[33]),
    .c(al_d6cb04b6[34]),
    .d(al_d6cb04b6[35]),
    .e(al_d6cb04b6[36]),
    .f(al_d6cb04b6[37]),
    .o(al_75ca1e75));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_e67818e8 (
    .a(al_b37de4b4),
    .b(al_7eb6704d),
    .c(al_d6cb04b6[44]),
    .d(al_d6cb04b6[45]),
    .e(al_d6cb04b6[50]),
    .f(al_d6cb04b6[51]),
    .o(al_4d58224c));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9166fb4b (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[23]),
    .d(al_96e7074d[0]),
    .o(al_3b7f0416[23]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3b2c95d0 (
    .a(al_d6cb04b6[40]),
    .b(al_d6cb04b6[41]),
    .c(al_d6cb04b6[42]),
    .d(al_d6cb04b6[43]),
    .o(al_f0189703));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_a6587af7 (
    .a(al_75ca1e75),
    .b(al_f0189703),
    .c(al_d6cb04b6[38]),
    .d(al_d6cb04b6[39]),
    .o(al_9fc9935f));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_d469bb84 (
    .a(al_d6cb04b6[52]),
    .b(al_d6cb04b6[53]),
    .c(al_d6cb04b6[54]),
    .d(al_96e7074d[9]),
    .o(al_b37de4b4));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_cf461ae3 (
    .a(al_d6cb04b6[46]),
    .b(al_d6cb04b6[47]),
    .c(al_d6cb04b6[48]),
    .d(al_d6cb04b6[49]),
    .o(al_7eb6704d));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_11c8b9b6 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[24]),
    .d(al_96e7074d[1]),
    .o(al_3b7f0416[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_be3161df (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[25]),
    .d(al_96e7074d[2]),
    .o(al_3b7f0416[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_7ce8b74 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[26]),
    .d(al_96e7074d[3]),
    .o(al_3b7f0416[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_18dbfceb (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[27]),
    .d(al_96e7074d[4]),
    .o(al_3b7f0416[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_b9d8be63 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[28]),
    .d(al_96e7074d[5]),
    .o(al_3b7f0416[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_8fb67e99 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[29]),
    .d(al_96e7074d[6]),
    .o(al_3b7f0416[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_889e55f4 (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[30]),
    .d(al_96e7074d[7]),
    .o(al_3b7f0416[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_9dacb12a (
    .a(al_9fc9935f),
    .b(al_4d58224c),
    .c(al_f7a9a92b[31]),
    .d(al_96e7074d[8]),
    .o(al_3b7f0416[31]));
  AL_DFF_X al_574b0a13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30922aac[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36d845bb[0]));
  AL_DFF_X al_39778347 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[22]));
  AL_DFF_X al_5858e220 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[23]));
  AL_DFF_X al_4667c1f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[24]));
  AL_DFF_X al_66c6deec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[25]));
  AL_DFF_X al_be577364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[26]));
  AL_DFF_X al_64f1e952 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[27]));
  AL_DFF_X al_1213b884 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[28]));
  AL_DFF_X al_dcc98efb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[29]));
  AL_DFF_X al_95380901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[30]));
  AL_DFF_X al_82457533 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[31]));
  AL_DFF_X al_f0ff413e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[32]));
  AL_DFF_X al_8f92702d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[33]));
  AL_DFF_X al_8be0a4d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[34]));
  AL_DFF_X al_e5e33e1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[35]));
  AL_DFF_X al_e7a6ff2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[36]));
  AL_DFF_X al_8e516f8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[37]));
  AL_DFF_X al_e66eb2b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[38]));
  AL_DFF_X al_b68c4f0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[39]));
  AL_DFF_X al_5b4abd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[40]));
  AL_DFF_X al_46d15407 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[41]));
  AL_DFF_X al_87f7d9e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[42]));
  AL_DFF_X al_acc51ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[43]));
  AL_DFF_X al_6830a2bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[44]));
  AL_DFF_X al_eded141d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[45]));
  AL_DFF_X al_144150ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[46]));
  AL_DFF_X al_2f0cc1cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[47]));
  AL_DFF_X al_9b9ec978 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[48]));
  AL_DFF_X al_eeff88d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[49]));
  AL_DFF_X al_1211bbf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[50]));
  AL_DFF_X al_1247c1f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[51]));
  AL_DFF_X al_c6053bee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[52]));
  AL_DFF_X al_d121c08f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[53]));
  AL_DFF_X al_dadcc19e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[8]));
  AL_DFF_X al_898f5520 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[9]));
  AL_DFF_X al_f61799d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[10]));
  AL_DFF_X al_63a42585 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[11]));
  AL_DFF_X al_6bd97037 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[12]));
  AL_DFF_X al_8afbb169 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[13]));
  AL_DFF_X al_51757c3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[14]));
  AL_DFF_X al_90a7f761 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[15]));
  AL_DFF_X al_fd77ea88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[16]));
  AL_DFF_X al_b9857e74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[17]));
  AL_DFF_X al_247320db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[0]));
  AL_DFF_X al_9ff3595 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[18]));
  AL_DFF_X al_9f18a690 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[19]));
  AL_DFF_X al_fa6e0364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[20]));
  AL_DFF_X al_1c5266d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[21]));
  AL_DFF_X al_37c6acc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[22]));
  AL_DFF_X al_13d9778 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[23]));
  AL_DFF_X al_7c0c3102 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[24]));
  AL_DFF_X al_76ef168c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[25]));
  AL_DFF_X al_8dcce430 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[26]));
  AL_DFF_X al_ffafa4bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[27]));
  AL_DFF_X al_cace1d7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[1]));
  AL_DFF_X al_38a24123 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[28]));
  AL_DFF_X al_1f364b73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[29]));
  AL_DFF_X al_e89100d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[30]));
  AL_DFF_X al_23d29d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[31]));
  AL_DFF_X al_c1695578 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[2]));
  AL_DFF_X al_af4ccdd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[3]));
  AL_DFF_X al_cb0090f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[4]));
  AL_DFF_X al_853a8f2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[5]));
  AL_DFF_X al_bfdaced4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[6]));
  AL_DFF_X al_47d7a0d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[7]));
  AL_DFF_X al_cfcf671f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[8]));
  AL_DFF_X al_a09f5853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d150e9d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[0]));
  AL_DFF_X al_17bc6b86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[1]));
  AL_DFF_X al_adc9fa19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[2]));
  AL_DFF_X al_5c0b6bfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[3]));
  AL_DFF_X al_a029932f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[4]));
  AL_DFF_X al_3641b87a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[5]));
  AL_DFF_X al_40b7a445 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[6]));
  AL_DFF_X al_c0e10d9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_fa2d4603 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .o(al_f058aa98));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1bfa61bf (
    .a(1'b0),
    .o({al_be714bda,open_n156}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_364d4d1c (
    .a(al_5283b07c[22]),
    .b(al_c1960abd[22]),
    .c(al_be714bda),
    .o({al_62b2844e,al_c855b680[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b596eab (
    .a(al_5283b07c[23]),
    .b(al_c1960abd[23]),
    .c(al_62b2844e),
    .o({al_23344b64,al_c855b680[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8e142b70 (
    .a(al_5283b07c[24]),
    .b(al_c1960abd[24]),
    .c(al_23344b64),
    .o({al_aa529150,al_c855b680[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_da020f26 (
    .a(al_5283b07c[25]),
    .b(al_c1960abd[25]),
    .c(al_aa529150),
    .o({al_d6b6abb7,al_c855b680[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2dc418bb (
    .a(al_5283b07c[26]),
    .b(al_c1960abd[26]),
    .c(al_d6b6abb7),
    .o({al_7cd30609,al_c855b680[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55832e89 (
    .a(al_5283b07c[27]),
    .b(al_c1960abd[27]),
    .c(al_7cd30609),
    .o({al_9765a29c,al_c855b680[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b36aedd6 (
    .a(al_5283b07c[28]),
    .b(al_c1960abd[28]),
    .c(al_9765a29c),
    .o({al_9d15fc0c,al_c855b680[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4e41d4c0 (
    .a(al_5283b07c[29]),
    .b(al_c1960abd[29]),
    .c(al_9d15fc0c),
    .o({al_8fcf5341,al_c855b680[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9ea535e (
    .a(al_5283b07c[30]),
    .b(al_c1960abd[30]),
    .c(al_8fcf5341),
    .o({al_5e79a92a,al_c855b680[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2b583e2 (
    .a(al_5283b07c[31]),
    .b(al_c1960abd[31]),
    .c(al_5e79a92a),
    .o({al_8fff10ae,al_c855b680[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d218d28 (
    .c(al_8fff10ae),
    .o({open_n159,al_c855b680[10]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_cbd377e5 (
    .a(al_c1960abd[42]),
    .b(al_c1960abd[43]),
    .c(al_c1960abd[44]),
    .d(al_c1960abd[45]),
    .e(al_c1960abd[46]),
    .f(al_c1960abd[47]),
    .o(al_bf66278b));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_b65429e1 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[22]),
    .e(al_c855b680[0]),
    .o(al_bcaebe78[22]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_ef71fb84 (
    .a(al_c1960abd[50]),
    .b(al_c1960abd[51]),
    .c(al_c1960abd[52]),
    .d(al_c1960abd[53]),
    .o(al_ec79a3f9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_e917d561 (
    .a(al_bf66278b),
    .b(al_ec79a3f9),
    .c(al_c1960abd[48]),
    .d(al_c1960abd[49]),
    .o(al_b02d6cd0));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_31488a58 (
    .a(al_c1960abd[36]),
    .b(al_c1960abd[37]),
    .c(al_c1960abd[38]),
    .d(al_c1960abd[39]),
    .e(al_c1960abd[40]),
    .f(al_c1960abd[41]),
    .o(al_c5e93959));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_b4bd6609 (
    .a(al_c1960abd[32]),
    .b(al_c1960abd[33]),
    .c(al_c1960abd[34]),
    .d(al_c1960abd[35]),
    .e(al_c855b680[10]),
    .o(al_dfb70c9));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_34e07716 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[23]),
    .e(al_c855b680[1]),
    .o(al_bcaebe78[23]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_56e3135 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[24]),
    .e(al_c855b680[2]),
    .o(al_bcaebe78[24]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_1cbd7002 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[25]),
    .e(al_c855b680[3]),
    .o(al_bcaebe78[25]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_672a66e0 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[26]),
    .e(al_c855b680[4]),
    .o(al_bcaebe78[26]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_60c80ba6 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[27]),
    .e(al_c855b680[5]),
    .o(al_bcaebe78[27]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_49c97c95 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[28]),
    .e(al_c855b680[6]),
    .o(al_bcaebe78[28]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_a0f6cea (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[29]),
    .e(al_c855b680[7]),
    .o(al_bcaebe78[29]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_bd1de708 (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[30]),
    .e(al_c855b680[8]),
    .o(al_bcaebe78[30]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((C*B*A))+D*E*~((C*B*A))+~(D)*E*(C*B*A)+D*E*(C*B*A))"),
    .INIT(32'hff807f00))
    al_1df0ccbb (
    .a(al_b02d6cd0),
    .b(al_c5e93959),
    .c(al_dfb70c9),
    .d(al_5283b07c[31]),
    .e(al_c855b680[9]),
    .o(al_bcaebe78[31]));
  AL_DFF_X al_c90585d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_36d845bb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b6a4daa[0]));
  AL_DFF_X al_e4a574bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[21]));
  AL_DFF_X al_39b55bf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[22]));
  AL_DFF_X al_11cc02bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[23]));
  AL_DFF_X al_804fbb51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[24]));
  AL_DFF_X al_dff05ff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[25]));
  AL_DFF_X al_e9932999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[26]));
  AL_DFF_X al_b4ad5d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[27]));
  AL_DFF_X al_9c21d93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[28]));
  AL_DFF_X al_2058bfee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[29]));
  AL_DFF_X al_61430c80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[30]));
  AL_DFF_X al_a1de8d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[31]));
  AL_DFF_X al_d26c59ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[32]));
  AL_DFF_X al_8309716f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[33]));
  AL_DFF_X al_4eb5bb4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[34]));
  AL_DFF_X al_168551a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[35]));
  AL_DFF_X al_b11d296f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[36]));
  AL_DFF_X al_b46c4d45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[37]));
  AL_DFF_X al_af58a36b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[38]));
  AL_DFF_X al_fd9a7217 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[39]));
  AL_DFF_X al_3049c75b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[40]));
  AL_DFF_X al_81434ad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[41]));
  AL_DFF_X al_82db834d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[42]));
  AL_DFF_X al_fdebac94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[43]));
  AL_DFF_X al_10c65464 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[44]));
  AL_DFF_X al_8cc78ffd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[45]));
  AL_DFF_X al_5653f9be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[46]));
  AL_DFF_X al_df9e6a5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[47]));
  AL_DFF_X al_25d9ab30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[48]));
  AL_DFF_X al_7f6149c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[49]));
  AL_DFF_X al_cf92fe55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[50]));
  AL_DFF_X al_f072bf1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[51]));
  AL_DFF_X al_fafa4f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[52]));
  AL_DFF_X al_e5c0deef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[8]));
  AL_DFF_X al_e69fce09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[9]));
  AL_DFF_X al_5945eb57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[10]));
  AL_DFF_X al_94973e49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[11]));
  AL_DFF_X al_b8c79f80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[12]));
  AL_DFF_X al_8ef49b3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[13]));
  AL_DFF_X al_26e0a8bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[14]));
  AL_DFF_X al_f0489817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[15]));
  AL_DFF_X al_42f4ad45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[16]));
  AL_DFF_X al_8c630f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[17]));
  AL_DFF_X al_3294900d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[0]));
  AL_DFF_X al_2332562b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[18]));
  AL_DFF_X al_80d3f8f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[19]));
  AL_DFF_X al_cfbe8dc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[20]));
  AL_DFF_X al_e3903be4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[21]));
  AL_DFF_X al_7a96ee43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[22]));
  AL_DFF_X al_a9d8dd44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[23]));
  AL_DFF_X al_771ddbe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[24]));
  AL_DFF_X al_303b2911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[25]));
  AL_DFF_X al_8a161fa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[26]));
  AL_DFF_X al_f5ed024e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[27]));
  AL_DFF_X al_7450b45d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[1]));
  AL_DFF_X al_942c503a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[28]));
  AL_DFF_X al_6670f26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[29]));
  AL_DFF_X al_fae1eb50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[30]));
  AL_DFF_X al_61d2ca3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[31]));
  AL_DFF_X al_310a5434 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[2]));
  AL_DFF_X al_a180323b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[3]));
  AL_DFF_X al_e361a27e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[4]));
  AL_DFF_X al_1dd11f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[5]));
  AL_DFF_X al_661bb2de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[6]));
  AL_DFF_X al_c5d4bfab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[7]));
  AL_DFF_X al_8b4c00b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[8]));
  AL_DFF_X al_9144a051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[9]));
  AL_DFF_X al_69edaf96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f058aa98),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[0]));
  AL_DFF_X al_95087f4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[1]));
  AL_DFF_X al_1837ab2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[2]));
  AL_DFF_X al_e5a7272c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[3]));
  AL_DFF_X al_2745e54d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[4]));
  AL_DFF_X al_5dd10ba1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[5]));
  AL_DFF_X al_b9bb8a3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[6]));
  AL_DFF_X al_6735a1a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[7]));
  AL_DFF_X al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ae5d831a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_DFF_X al_65d1adb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[31]));
  AL_DFF_X al_f66a344 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[32]));
  AL_DFF_X al_f617f18d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[33]));
  AL_DFF_X al_9faa4a4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[34]));
  AL_DFF_X al_fc166c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[35]));
  AL_DFF_X al_4c8ce131 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[36]));
  AL_DFF_X al_2637942e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[37]));
  AL_DFF_X al_a7daa706 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[38]));
  AL_DFF_X al_a3b5c5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[39]));
  AL_DFF_X al_9ec017c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[40]));
  AL_DFF_X al_61f52352 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[41]));
  AL_DFF_X al_3e920ff5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[42]));
  AL_DFF_X al_c2e2478e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[43]));
  AL_DFF_X al_8eba0e17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[44]));
  AL_DFF_X al_5c5b7a6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[45]));
  AL_DFF_X al_523a6904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[46]));
  AL_DFF_X al_7ac71266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[47]));
  AL_DFF_X al_138d45d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[48]));
  AL_DFF_X al_fde31f80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[49]));
  AL_DFF_X al_bd637999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[50]));
  AL_DFF_X al_cda6c19b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[51]));
  AL_DFF_X al_abb9599d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[52]));
  AL_DFF_X al_8de7e0a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[53]));
  AL_DFF_X al_1fe8680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[54]));
  AL_DFF_X al_92a923a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[55]));
  AL_DFF_X al_5a3580e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[56]));
  AL_DFF_X al_7ac7438a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[57]));
  AL_DFF_X al_48b78abc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[58]));
  AL_DFF_X al_40261b07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[59]));
  AL_DFF_X al_7b4b93f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[60]));
  AL_DFF_X al_97ffc327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[61]));
  AL_DFF_X al_a8743118 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[62]));
  AL_DFF_X al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[8]));
  AL_DFF_X al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[9]));
  AL_DFF_X al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[10]));
  AL_DFF_X al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[11]));
  AL_DFF_X al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[12]));
  AL_DFF_X al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[13]));
  AL_DFF_X al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[14]));
  AL_DFF_X al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[15]));
  AL_DFF_X al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[16]));
  AL_DFF_X al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[17]));
  AL_DFF_X al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[0]));
  AL_DFF_X al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[18]));
  AL_DFF_X al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[19]));
  AL_DFF_X al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[20]));
  AL_DFF_X al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[21]));
  AL_DFF_X al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[22]));
  AL_DFF_X al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[23]));
  AL_DFF_X al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[24]));
  AL_DFF_X al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[25]));
  AL_DFF_X al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[26]));
  AL_DFF_X al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[27]));
  AL_DFF_X al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[1]));
  AL_DFF_X al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[28]));
  AL_DFF_X al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[29]));
  AL_DFF_X al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[30]));
  AL_DFF_X al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[31]));
  AL_DFF_X al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[2]));
  AL_DFF_X al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[3]));
  AL_DFF_X al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[4]));
  AL_DFF_X al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[5]));
  AL_DFF_X al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[6]));
  AL_DFF_X al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[7]));
  AL_DFF_X al_596b0fc4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_X al_5cfa2c1e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_X al_c56c02f8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_X al_60ec2662 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_X al_ea3f598e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_X al_dd4ae85d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_X al_e2aa8055 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_X al_82aa8ce (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_X al_7f911c70 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_X al_8908ba38 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_X al_16ad90bc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_X al_2149b062 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_X al_56d82898 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_X al_c8bec57f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_X al_1f071837 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_X al_9acbb644 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_X al_286bd0de (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_X al_7e8bb9f7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_X al_d4e324dc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_X al_bcaf406d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_X al_20d194ca (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[27]));
  AL_DFF_X al_e1044ec0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_X al_6402198 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[28]));
  AL_DFF_X al_3f7239b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[29]));
  AL_DFF_X al_33cd891 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[30]));
  AL_DFF_X al_28b9e853 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[31]));
  AL_DFF_X al_16da6de4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_X al_e819e904 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_X al_4990808d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_X al_d51e17ed (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_X al_b67f884b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_X al_ff3308ea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_18157fe8[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_X al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_X al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_X al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_X al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_X al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_X al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_X al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_X al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_X al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_X al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_X al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_X al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_X al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_X al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_X al_c179532 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[21]));
  AL_DFF_X al_7d105784 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[22]));
  AL_DFF_X al_573a0a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[23]));
  AL_DFF_X al_d0deffcb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[24]));
  AL_DFF_X al_150254f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[25]));
  AL_DFF_X al_47f1ba67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[26]));
  AL_DFF_X al_3f6c28d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[27]));
  AL_DFF_X al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_X al_930b6560 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[28]));
  AL_DFF_X al_46a886ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[29]));
  AL_DFF_X al_5c18d1b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[30]));
  AL_DFF_X al_f94ac09a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[31]));
  AL_DFF_X al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_X al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_X al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_X al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_X al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_X al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3519ff8d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_DFF_X al_f6de6753 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(start),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51794c84));

endmodule 

